# ________________________________________________________________________________________________
# 
# 
#             Synchronous RVT Periphery One-Port Register File Compiler
# 
#                 UMC 55nm Low K Low Power Logic Process
# 
# ________________________________________________________________________________________________
# 
#               
#         Copyright (C) 2020 Faraday Technology Corporation. All Rights Reserved.       
#                
#         This source code is an unpublished work belongs to Faraday Technology Corporation       
#         It is considered a trade secret and is not to be divulged or       
#         used by parties who have not received written authorization from       
#         Faraday Technology Corporation       
#                
#         Faraday's home page can be found at: http://www.faraday-tech.com/       
#                
# ________________________________________________________________________________________________
# 
#        IP Name            :  FSF0L_A_SY                                    
#        IP Version         :  1.5.0                                         
#        IP Release Status  :  Active                                        
#        Word               :  512                                           
#        Bit                :  32                                            
#        Byte               :  4                                             
#        Mux                :  2                                             
#        Output Loading     :  0.01                                          
#        Clock Input Slew   :  0.008                                         
#        Data Input Slew    :  0.008                                         
#        Ring Type          :  Ring Shape Model                              
#        Ring Layer         :  2233                                          
#        Ring Width         :  2                                             
#        Bus Format         :  1                                             
#        Memaker Path       :  /workspace/technology/umc/55nm_201908/memlib  
#        GUI Version        :  m20130120                                     
#        Date               :  2020/07/14 13:57:08                           
# ________________________________________________________________________________________________
# 

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
MACRO SYLA55_512X32X4CM2
CLASS BLOCK ;
FOREIGN SYLA55_512X32X4CM2 0.000 0.000 ;
ORIGIN 0.000 0.000 ;
SIZE 298.405 BY 164.840 ;
SYMMETRY x y r90 ;
SITE core ;
PIN DI[63]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 138.315 4.600 138.475 4.700 ;
  LAYER ME2 ;
  RECT 138.315 4.600 138.475 4.700 ;
  LAYER ME1 ;
  RECT 138.315 4.600 138.475 4.700 ;
  LAYER VI1 ;
  RECT 138.345 4.600 138.445 4.700 ;
  LAYER VI2 ;
  RECT 138.345 4.600 138.445 4.700 ;
  LAYER VI3 ;
  RECT 138.345 4.600 138.445 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[63]
PIN DO[63]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 139.715 4.600 139.875 4.700 ;
  LAYER ME2 ;
  RECT 139.715 4.600 139.875 4.700 ;
  LAYER ME1 ;
  RECT 139.715 4.600 139.875 4.700 ;
  LAYER VI1 ;
  RECT 139.745 4.600 139.845 4.700 ;
  LAYER VI2 ;
  RECT 139.745 4.600 139.845 4.700 ;
  LAYER VI3 ;
  RECT 139.745 4.600 139.845 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[63]
PIN DI[62]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 136.215 4.600 136.375 4.700 ;
  LAYER ME2 ;
  RECT 136.215 4.600 136.375 4.700 ;
  LAYER ME1 ;
  RECT 136.215 4.600 136.375 4.700 ;
  LAYER VI1 ;
  RECT 136.245 4.600 136.345 4.700 ;
  LAYER VI2 ;
  RECT 136.245 4.600 136.345 4.700 ;
  LAYER VI3 ;
  RECT 136.245 4.600 136.345 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[62]
PIN DO[62]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 137.615 4.600 137.775 4.700 ;
  LAYER ME2 ;
  RECT 137.615 4.600 137.775 4.700 ;
  LAYER ME1 ;
  RECT 137.615 4.600 137.775 4.700 ;
  LAYER VI1 ;
  RECT 137.645 4.600 137.745 4.700 ;
  LAYER VI2 ;
  RECT 137.645 4.600 137.745 4.700 ;
  LAYER VI3 ;
  RECT 137.645 4.600 137.745 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[62]
PIN DI[61]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 134.115 4.600 134.275 4.700 ;
  LAYER ME2 ;
  RECT 134.115 4.600 134.275 4.700 ;
  LAYER ME1 ;
  RECT 134.115 4.600 134.275 4.700 ;
  LAYER VI1 ;
  RECT 134.145 4.600 134.245 4.700 ;
  LAYER VI2 ;
  RECT 134.145 4.600 134.245 4.700 ;
  LAYER VI3 ;
  RECT 134.145 4.600 134.245 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[61]
PIN DO[61]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 135.515 4.600 135.675 4.700 ;
  LAYER ME2 ;
  RECT 135.515 4.600 135.675 4.700 ;
  LAYER ME1 ;
  RECT 135.515 4.600 135.675 4.700 ;
  LAYER VI1 ;
  RECT 135.545 4.600 135.645 4.700 ;
  LAYER VI2 ;
  RECT 135.545 4.600 135.645 4.700 ;
  LAYER VI3 ;
  RECT 135.545 4.600 135.645 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[61]
PIN DI[60]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 132.015 4.600 132.175 4.700 ;
  LAYER ME2 ;
  RECT 132.015 4.600 132.175 4.700 ;
  LAYER ME1 ;
  RECT 132.015 4.600 132.175 4.700 ;
  LAYER VI1 ;
  RECT 132.045 4.600 132.145 4.700 ;
  LAYER VI2 ;
  RECT 132.045 4.600 132.145 4.700 ;
  LAYER VI3 ;
  RECT 132.045 4.600 132.145 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[60]
PIN DO[60]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 133.415 4.600 133.575 4.700 ;
  LAYER ME2 ;
  RECT 133.415 4.600 133.575 4.700 ;
  LAYER ME1 ;
  RECT 133.415 4.600 133.575 4.700 ;
  LAYER VI1 ;
  RECT 133.445 4.600 133.545 4.700 ;
  LAYER VI2 ;
  RECT 133.445 4.600 133.545 4.700 ;
  LAYER VI3 ;
  RECT 133.445 4.600 133.545 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[60]
PIN DI[59]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 129.915 4.600 130.075 4.700 ;
  LAYER ME2 ;
  RECT 129.915 4.600 130.075 4.700 ;
  LAYER ME1 ;
  RECT 129.915 4.600 130.075 4.700 ;
  LAYER VI1 ;
  RECT 129.945 4.600 130.045 4.700 ;
  LAYER VI2 ;
  RECT 129.945 4.600 130.045 4.700 ;
  LAYER VI3 ;
  RECT 129.945 4.600 130.045 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[59]
PIN DO[59]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 131.315 4.600 131.475 4.700 ;
  LAYER ME2 ;
  RECT 131.315 4.600 131.475 4.700 ;
  LAYER ME1 ;
  RECT 131.315 4.600 131.475 4.700 ;
  LAYER VI1 ;
  RECT 131.345 4.600 131.445 4.700 ;
  LAYER VI2 ;
  RECT 131.345 4.600 131.445 4.700 ;
  LAYER VI3 ;
  RECT 131.345 4.600 131.445 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[59]
PIN DI[58]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 127.815 4.600 127.975 4.700 ;
  LAYER ME2 ;
  RECT 127.815 4.600 127.975 4.700 ;
  LAYER ME1 ;
  RECT 127.815 4.600 127.975 4.700 ;
  LAYER VI1 ;
  RECT 127.845 4.600 127.945 4.700 ;
  LAYER VI2 ;
  RECT 127.845 4.600 127.945 4.700 ;
  LAYER VI3 ;
  RECT 127.845 4.600 127.945 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[58]
PIN DO[58]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 129.215 4.600 129.375 4.700 ;
  LAYER ME2 ;
  RECT 129.215 4.600 129.375 4.700 ;
  LAYER ME1 ;
  RECT 129.215 4.600 129.375 4.700 ;
  LAYER VI1 ;
  RECT 129.245 4.600 129.345 4.700 ;
  LAYER VI2 ;
  RECT 129.245 4.600 129.345 4.700 ;
  LAYER VI3 ;
  RECT 129.245 4.600 129.345 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[58]
PIN DI[57]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 125.715 4.600 125.875 4.700 ;
  LAYER ME2 ;
  RECT 125.715 4.600 125.875 4.700 ;
  LAYER ME1 ;
  RECT 125.715 4.600 125.875 4.700 ;
  LAYER VI1 ;
  RECT 125.745 4.600 125.845 4.700 ;
  LAYER VI2 ;
  RECT 125.745 4.600 125.845 4.700 ;
  LAYER VI3 ;
  RECT 125.745 4.600 125.845 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[57]
PIN DO[57]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 127.115 4.600 127.275 4.700 ;
  LAYER ME2 ;
  RECT 127.115 4.600 127.275 4.700 ;
  LAYER ME1 ;
  RECT 127.115 4.600 127.275 4.700 ;
  LAYER VI1 ;
  RECT 127.145 4.600 127.245 4.700 ;
  LAYER VI2 ;
  RECT 127.145 4.600 127.245 4.700 ;
  LAYER VI3 ;
  RECT 127.145 4.600 127.245 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[57]
PIN DI[56]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 123.615 4.600 123.775 4.700 ;
  LAYER ME2 ;
  RECT 123.615 4.600 123.775 4.700 ;
  LAYER ME1 ;
  RECT 123.615 4.600 123.775 4.700 ;
  LAYER VI1 ;
  RECT 123.645 4.600 123.745 4.700 ;
  LAYER VI2 ;
  RECT 123.645 4.600 123.745 4.700 ;
  LAYER VI3 ;
  RECT 123.645 4.600 123.745 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[56]
PIN DO[56]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 125.015 4.600 125.175 4.700 ;
  LAYER ME2 ;
  RECT 125.015 4.600 125.175 4.700 ;
  LAYER ME1 ;
  RECT 125.015 4.600 125.175 4.700 ;
  LAYER VI1 ;
  RECT 125.045 4.600 125.145 4.700 ;
  LAYER VI2 ;
  RECT 125.045 4.600 125.145 4.700 ;
  LAYER VI3 ;
  RECT 125.045 4.600 125.145 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[56]
PIN DI[55]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 121.515 4.600 121.675 4.700 ;
  LAYER ME2 ;
  RECT 121.515 4.600 121.675 4.700 ;
  LAYER ME1 ;
  RECT 121.515 4.600 121.675 4.700 ;
  LAYER VI1 ;
  RECT 121.545 4.600 121.645 4.700 ;
  LAYER VI2 ;
  RECT 121.545 4.600 121.645 4.700 ;
  LAYER VI3 ;
  RECT 121.545 4.600 121.645 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[55]
PIN DO[55]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 122.915 4.600 123.075 4.700 ;
  LAYER ME2 ;
  RECT 122.915 4.600 123.075 4.700 ;
  LAYER ME1 ;
  RECT 122.915 4.600 123.075 4.700 ;
  LAYER VI1 ;
  RECT 122.945 4.600 123.045 4.700 ;
  LAYER VI2 ;
  RECT 122.945 4.600 123.045 4.700 ;
  LAYER VI3 ;
  RECT 122.945 4.600 123.045 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[55]
PIN DI[54]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 119.415 4.600 119.575 4.700 ;
  LAYER ME2 ;
  RECT 119.415 4.600 119.575 4.700 ;
  LAYER ME1 ;
  RECT 119.415 4.600 119.575 4.700 ;
  LAYER VI1 ;
  RECT 119.445 4.600 119.545 4.700 ;
  LAYER VI2 ;
  RECT 119.445 4.600 119.545 4.700 ;
  LAYER VI3 ;
  RECT 119.445 4.600 119.545 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[54]
PIN DO[54]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 120.815 4.600 120.975 4.700 ;
  LAYER ME2 ;
  RECT 120.815 4.600 120.975 4.700 ;
  LAYER ME1 ;
  RECT 120.815 4.600 120.975 4.700 ;
  LAYER VI1 ;
  RECT 120.845 4.600 120.945 4.700 ;
  LAYER VI2 ;
  RECT 120.845 4.600 120.945 4.700 ;
  LAYER VI3 ;
  RECT 120.845 4.600 120.945 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[54]
PIN DI[53]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 117.315 4.600 117.475 4.700 ;
  LAYER ME2 ;
  RECT 117.315 4.600 117.475 4.700 ;
  LAYER ME1 ;
  RECT 117.315 4.600 117.475 4.700 ;
  LAYER VI1 ;
  RECT 117.345 4.600 117.445 4.700 ;
  LAYER VI2 ;
  RECT 117.345 4.600 117.445 4.700 ;
  LAYER VI3 ;
  RECT 117.345 4.600 117.445 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[53]
PIN DO[53]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 118.715 4.600 118.875 4.700 ;
  LAYER ME2 ;
  RECT 118.715 4.600 118.875 4.700 ;
  LAYER ME1 ;
  RECT 118.715 4.600 118.875 4.700 ;
  LAYER VI1 ;
  RECT 118.745 4.600 118.845 4.700 ;
  LAYER VI2 ;
  RECT 118.745 4.600 118.845 4.700 ;
  LAYER VI3 ;
  RECT 118.745 4.600 118.845 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[53]
PIN DI[52]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 115.215 4.600 115.375 4.700 ;
  LAYER ME2 ;
  RECT 115.215 4.600 115.375 4.700 ;
  LAYER ME1 ;
  RECT 115.215 4.600 115.375 4.700 ;
  LAYER VI1 ;
  RECT 115.245 4.600 115.345 4.700 ;
  LAYER VI2 ;
  RECT 115.245 4.600 115.345 4.700 ;
  LAYER VI3 ;
  RECT 115.245 4.600 115.345 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[52]
PIN DO[52]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 116.615 4.600 116.775 4.700 ;
  LAYER ME2 ;
  RECT 116.615 4.600 116.775 4.700 ;
  LAYER ME1 ;
  RECT 116.615 4.600 116.775 4.700 ;
  LAYER VI1 ;
  RECT 116.645 4.600 116.745 4.700 ;
  LAYER VI2 ;
  RECT 116.645 4.600 116.745 4.700 ;
  LAYER VI3 ;
  RECT 116.645 4.600 116.745 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[52]
PIN DI[51]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 113.115 4.600 113.275 4.700 ;
  LAYER ME2 ;
  RECT 113.115 4.600 113.275 4.700 ;
  LAYER ME1 ;
  RECT 113.115 4.600 113.275 4.700 ;
  LAYER VI1 ;
  RECT 113.145 4.600 113.245 4.700 ;
  LAYER VI2 ;
  RECT 113.145 4.600 113.245 4.700 ;
  LAYER VI3 ;
  RECT 113.145 4.600 113.245 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[51]
PIN DO[51]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 114.515 4.600 114.675 4.700 ;
  LAYER ME2 ;
  RECT 114.515 4.600 114.675 4.700 ;
  LAYER ME1 ;
  RECT 114.515 4.600 114.675 4.700 ;
  LAYER VI1 ;
  RECT 114.545 4.600 114.645 4.700 ;
  LAYER VI2 ;
  RECT 114.545 4.600 114.645 4.700 ;
  LAYER VI3 ;
  RECT 114.545 4.600 114.645 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[51]
PIN DI[50]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 111.015 4.600 111.175 4.700 ;
  LAYER ME2 ;
  RECT 111.015 4.600 111.175 4.700 ;
  LAYER ME1 ;
  RECT 111.015 4.600 111.175 4.700 ;
  LAYER VI1 ;
  RECT 111.045 4.600 111.145 4.700 ;
  LAYER VI2 ;
  RECT 111.045 4.600 111.145 4.700 ;
  LAYER VI3 ;
  RECT 111.045 4.600 111.145 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[50]
PIN DO[50]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 112.415 4.600 112.575 4.700 ;
  LAYER ME2 ;
  RECT 112.415 4.600 112.575 4.700 ;
  LAYER ME1 ;
  RECT 112.415 4.600 112.575 4.700 ;
  LAYER VI1 ;
  RECT 112.445 4.600 112.545 4.700 ;
  LAYER VI2 ;
  RECT 112.445 4.600 112.545 4.700 ;
  LAYER VI3 ;
  RECT 112.445 4.600 112.545 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[50]
PIN DI[49]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 108.915 4.600 109.075 4.700 ;
  LAYER ME2 ;
  RECT 108.915 4.600 109.075 4.700 ;
  LAYER ME1 ;
  RECT 108.915 4.600 109.075 4.700 ;
  LAYER VI1 ;
  RECT 108.945 4.600 109.045 4.700 ;
  LAYER VI2 ;
  RECT 108.945 4.600 109.045 4.700 ;
  LAYER VI3 ;
  RECT 108.945 4.600 109.045 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[49]
PIN DO[49]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 110.315 4.600 110.475 4.700 ;
  LAYER ME2 ;
  RECT 110.315 4.600 110.475 4.700 ;
  LAYER ME1 ;
  RECT 110.315 4.600 110.475 4.700 ;
  LAYER VI1 ;
  RECT 110.345 4.600 110.445 4.700 ;
  LAYER VI2 ;
  RECT 110.345 4.600 110.445 4.700 ;
  LAYER VI3 ;
  RECT 110.345 4.600 110.445 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[49]
PIN DI[48]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 106.815 4.600 106.975 4.700 ;
  LAYER ME2 ;
  RECT 106.815 4.600 106.975 4.700 ;
  LAYER ME1 ;
  RECT 106.815 4.600 106.975 4.700 ;
  LAYER VI1 ;
  RECT 106.845 4.600 106.945 4.700 ;
  LAYER VI2 ;
  RECT 106.845 4.600 106.945 4.700 ;
  LAYER VI3 ;
  RECT 106.845 4.600 106.945 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[48]
PIN DO[48]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 108.215 4.600 108.375 4.700 ;
  LAYER ME2 ;
  RECT 108.215 4.600 108.375 4.700 ;
  LAYER ME1 ;
  RECT 108.215 4.600 108.375 4.700 ;
  LAYER VI1 ;
  RECT 108.245 4.600 108.345 4.700 ;
  LAYER VI2 ;
  RECT 108.245 4.600 108.345 4.700 ;
  LAYER VI3 ;
  RECT 108.245 4.600 108.345 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[48]
PIN DI[47]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 104.715 4.600 104.875 4.700 ;
  LAYER ME2 ;
  RECT 104.715 4.600 104.875 4.700 ;
  LAYER ME1 ;
  RECT 104.715 4.600 104.875 4.700 ;
  LAYER VI1 ;
  RECT 104.745 4.600 104.845 4.700 ;
  LAYER VI2 ;
  RECT 104.745 4.600 104.845 4.700 ;
  LAYER VI3 ;
  RECT 104.745 4.600 104.845 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[47]
PIN DO[47]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 106.115 4.600 106.275 4.700 ;
  LAYER ME2 ;
  RECT 106.115 4.600 106.275 4.700 ;
  LAYER ME1 ;
  RECT 106.115 4.600 106.275 4.700 ;
  LAYER VI1 ;
  RECT 106.145 4.600 106.245 4.700 ;
  LAYER VI2 ;
  RECT 106.145 4.600 106.245 4.700 ;
  LAYER VI3 ;
  RECT 106.145 4.600 106.245 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[47]
PIN DI[46]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 102.615 4.600 102.775 4.700 ;
  LAYER ME2 ;
  RECT 102.615 4.600 102.775 4.700 ;
  LAYER ME1 ;
  RECT 102.615 4.600 102.775 4.700 ;
  LAYER VI1 ;
  RECT 102.645 4.600 102.745 4.700 ;
  LAYER VI2 ;
  RECT 102.645 4.600 102.745 4.700 ;
  LAYER VI3 ;
  RECT 102.645 4.600 102.745 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[46]
PIN DO[46]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 104.015 4.600 104.175 4.700 ;
  LAYER ME2 ;
  RECT 104.015 4.600 104.175 4.700 ;
  LAYER ME1 ;
  RECT 104.015 4.600 104.175 4.700 ;
  LAYER VI1 ;
  RECT 104.045 4.600 104.145 4.700 ;
  LAYER VI2 ;
  RECT 104.045 4.600 104.145 4.700 ;
  LAYER VI3 ;
  RECT 104.045 4.600 104.145 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[46]
PIN DI[45]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 100.515 4.600 100.675 4.700 ;
  LAYER ME2 ;
  RECT 100.515 4.600 100.675 4.700 ;
  LAYER ME1 ;
  RECT 100.515 4.600 100.675 4.700 ;
  LAYER VI1 ;
  RECT 100.545 4.600 100.645 4.700 ;
  LAYER VI2 ;
  RECT 100.545 4.600 100.645 4.700 ;
  LAYER VI3 ;
  RECT 100.545 4.600 100.645 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[45]
PIN DO[45]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 101.915 4.600 102.075 4.700 ;
  LAYER ME2 ;
  RECT 101.915 4.600 102.075 4.700 ;
  LAYER ME1 ;
  RECT 101.915 4.600 102.075 4.700 ;
  LAYER VI1 ;
  RECT 101.945 4.600 102.045 4.700 ;
  LAYER VI2 ;
  RECT 101.945 4.600 102.045 4.700 ;
  LAYER VI3 ;
  RECT 101.945 4.600 102.045 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[45]
PIN DI[44]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 98.415 4.600 98.575 4.700 ;
  LAYER ME2 ;
  RECT 98.415 4.600 98.575 4.700 ;
  LAYER ME1 ;
  RECT 98.415 4.600 98.575 4.700 ;
  LAYER VI1 ;
  RECT 98.445 4.600 98.545 4.700 ;
  LAYER VI2 ;
  RECT 98.445 4.600 98.545 4.700 ;
  LAYER VI3 ;
  RECT 98.445 4.600 98.545 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[44]
PIN DO[44]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 99.815 4.600 99.975 4.700 ;
  LAYER ME2 ;
  RECT 99.815 4.600 99.975 4.700 ;
  LAYER ME1 ;
  RECT 99.815 4.600 99.975 4.700 ;
  LAYER VI1 ;
  RECT 99.845 4.600 99.945 4.700 ;
  LAYER VI2 ;
  RECT 99.845 4.600 99.945 4.700 ;
  LAYER VI3 ;
  RECT 99.845 4.600 99.945 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[44]
PIN DI[43]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 96.315 4.600 96.475 4.700 ;
  LAYER ME2 ;
  RECT 96.315 4.600 96.475 4.700 ;
  LAYER ME1 ;
  RECT 96.315 4.600 96.475 4.700 ;
  LAYER VI1 ;
  RECT 96.345 4.600 96.445 4.700 ;
  LAYER VI2 ;
  RECT 96.345 4.600 96.445 4.700 ;
  LAYER VI3 ;
  RECT 96.345 4.600 96.445 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[43]
PIN DO[43]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 97.715 4.600 97.875 4.700 ;
  LAYER ME2 ;
  RECT 97.715 4.600 97.875 4.700 ;
  LAYER ME1 ;
  RECT 97.715 4.600 97.875 4.700 ;
  LAYER VI1 ;
  RECT 97.745 4.600 97.845 4.700 ;
  LAYER VI2 ;
  RECT 97.745 4.600 97.845 4.700 ;
  LAYER VI3 ;
  RECT 97.745 4.600 97.845 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[43]
PIN DI[42]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 94.215 4.600 94.375 4.700 ;
  LAYER ME2 ;
  RECT 94.215 4.600 94.375 4.700 ;
  LAYER ME1 ;
  RECT 94.215 4.600 94.375 4.700 ;
  LAYER VI1 ;
  RECT 94.245 4.600 94.345 4.700 ;
  LAYER VI2 ;
  RECT 94.245 4.600 94.345 4.700 ;
  LAYER VI3 ;
  RECT 94.245 4.600 94.345 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[42]
PIN DO[42]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 95.615 4.600 95.775 4.700 ;
  LAYER ME2 ;
  RECT 95.615 4.600 95.775 4.700 ;
  LAYER ME1 ;
  RECT 95.615 4.600 95.775 4.700 ;
  LAYER VI1 ;
  RECT 95.645 4.600 95.745 4.700 ;
  LAYER VI2 ;
  RECT 95.645 4.600 95.745 4.700 ;
  LAYER VI3 ;
  RECT 95.645 4.600 95.745 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[42]
PIN DI[41]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 92.115 4.600 92.275 4.700 ;
  LAYER ME2 ;
  RECT 92.115 4.600 92.275 4.700 ;
  LAYER ME1 ;
  RECT 92.115 4.600 92.275 4.700 ;
  LAYER VI1 ;
  RECT 92.145 4.600 92.245 4.700 ;
  LAYER VI2 ;
  RECT 92.145 4.600 92.245 4.700 ;
  LAYER VI3 ;
  RECT 92.145 4.600 92.245 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[41]
PIN DO[41]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 93.515 4.600 93.675 4.700 ;
  LAYER ME2 ;
  RECT 93.515 4.600 93.675 4.700 ;
  LAYER ME1 ;
  RECT 93.515 4.600 93.675 4.700 ;
  LAYER VI1 ;
  RECT 93.545 4.600 93.645 4.700 ;
  LAYER VI2 ;
  RECT 93.545 4.600 93.645 4.700 ;
  LAYER VI3 ;
  RECT 93.545 4.600 93.645 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[41]
PIN DI[40]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 90.015 4.600 90.175 4.700 ;
  LAYER ME2 ;
  RECT 90.015 4.600 90.175 4.700 ;
  LAYER ME1 ;
  RECT 90.015 4.600 90.175 4.700 ;
  LAYER VI1 ;
  RECT 90.045 4.600 90.145 4.700 ;
  LAYER VI2 ;
  RECT 90.045 4.600 90.145 4.700 ;
  LAYER VI3 ;
  RECT 90.045 4.600 90.145 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[40]
PIN DO[40]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 91.415 4.600 91.575 4.700 ;
  LAYER ME2 ;
  RECT 91.415 4.600 91.575 4.700 ;
  LAYER ME1 ;
  RECT 91.415 4.600 91.575 4.700 ;
  LAYER VI1 ;
  RECT 91.445 4.600 91.545 4.700 ;
  LAYER VI2 ;
  RECT 91.445 4.600 91.545 4.700 ;
  LAYER VI3 ;
  RECT 91.445 4.600 91.545 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[40]
PIN DI[39]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 87.915 4.600 88.075 4.700 ;
  LAYER ME2 ;
  RECT 87.915 4.600 88.075 4.700 ;
  LAYER ME1 ;
  RECT 87.915 4.600 88.075 4.700 ;
  LAYER VI1 ;
  RECT 87.945 4.600 88.045 4.700 ;
  LAYER VI2 ;
  RECT 87.945 4.600 88.045 4.700 ;
  LAYER VI3 ;
  RECT 87.945 4.600 88.045 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[39]
PIN DO[39]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 89.315 4.600 89.475 4.700 ;
  LAYER ME2 ;
  RECT 89.315 4.600 89.475 4.700 ;
  LAYER ME1 ;
  RECT 89.315 4.600 89.475 4.700 ;
  LAYER VI1 ;
  RECT 89.345 4.600 89.445 4.700 ;
  LAYER VI2 ;
  RECT 89.345 4.600 89.445 4.700 ;
  LAYER VI3 ;
  RECT 89.345 4.600 89.445 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[39]
PIN DI[38]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 85.815 4.600 85.975 4.700 ;
  LAYER ME2 ;
  RECT 85.815 4.600 85.975 4.700 ;
  LAYER ME1 ;
  RECT 85.815 4.600 85.975 4.700 ;
  LAYER VI1 ;
  RECT 85.845 4.600 85.945 4.700 ;
  LAYER VI2 ;
  RECT 85.845 4.600 85.945 4.700 ;
  LAYER VI3 ;
  RECT 85.845 4.600 85.945 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[38]
PIN DO[38]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 87.215 4.600 87.375 4.700 ;
  LAYER ME2 ;
  RECT 87.215 4.600 87.375 4.700 ;
  LAYER ME1 ;
  RECT 87.215 4.600 87.375 4.700 ;
  LAYER VI1 ;
  RECT 87.245 4.600 87.345 4.700 ;
  LAYER VI2 ;
  RECT 87.245 4.600 87.345 4.700 ;
  LAYER VI3 ;
  RECT 87.245 4.600 87.345 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[38]
PIN DI[37]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 83.715 4.600 83.875 4.700 ;
  LAYER ME2 ;
  RECT 83.715 4.600 83.875 4.700 ;
  LAYER ME1 ;
  RECT 83.715 4.600 83.875 4.700 ;
  LAYER VI1 ;
  RECT 83.745 4.600 83.845 4.700 ;
  LAYER VI2 ;
  RECT 83.745 4.600 83.845 4.700 ;
  LAYER VI3 ;
  RECT 83.745 4.600 83.845 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[37]
PIN DO[37]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 85.115 4.600 85.275 4.700 ;
  LAYER ME2 ;
  RECT 85.115 4.600 85.275 4.700 ;
  LAYER ME1 ;
  RECT 85.115 4.600 85.275 4.700 ;
  LAYER VI1 ;
  RECT 85.145 4.600 85.245 4.700 ;
  LAYER VI2 ;
  RECT 85.145 4.600 85.245 4.700 ;
  LAYER VI3 ;
  RECT 85.145 4.600 85.245 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[37]
PIN DI[36]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 81.615 4.600 81.775 4.700 ;
  LAYER ME2 ;
  RECT 81.615 4.600 81.775 4.700 ;
  LAYER ME1 ;
  RECT 81.615 4.600 81.775 4.700 ;
  LAYER VI1 ;
  RECT 81.645 4.600 81.745 4.700 ;
  LAYER VI2 ;
  RECT 81.645 4.600 81.745 4.700 ;
  LAYER VI3 ;
  RECT 81.645 4.600 81.745 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[36]
PIN DO[36]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 83.015 4.600 83.175 4.700 ;
  LAYER ME2 ;
  RECT 83.015 4.600 83.175 4.700 ;
  LAYER ME1 ;
  RECT 83.015 4.600 83.175 4.700 ;
  LAYER VI1 ;
  RECT 83.045 4.600 83.145 4.700 ;
  LAYER VI2 ;
  RECT 83.045 4.600 83.145 4.700 ;
  LAYER VI3 ;
  RECT 83.045 4.600 83.145 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[36]
PIN DI[35]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 79.515 4.600 79.675 4.700 ;
  LAYER ME2 ;
  RECT 79.515 4.600 79.675 4.700 ;
  LAYER ME1 ;
  RECT 79.515 4.600 79.675 4.700 ;
  LAYER VI1 ;
  RECT 79.545 4.600 79.645 4.700 ;
  LAYER VI2 ;
  RECT 79.545 4.600 79.645 4.700 ;
  LAYER VI3 ;
  RECT 79.545 4.600 79.645 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[35]
PIN DO[35]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 80.915 4.600 81.075 4.700 ;
  LAYER ME2 ;
  RECT 80.915 4.600 81.075 4.700 ;
  LAYER ME1 ;
  RECT 80.915 4.600 81.075 4.700 ;
  LAYER VI1 ;
  RECT 80.945 4.600 81.045 4.700 ;
  LAYER VI2 ;
  RECT 80.945 4.600 81.045 4.700 ;
  LAYER VI3 ;
  RECT 80.945 4.600 81.045 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[35]
PIN DI[34]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 77.415 4.600 77.575 4.700 ;
  LAYER ME2 ;
  RECT 77.415 4.600 77.575 4.700 ;
  LAYER ME1 ;
  RECT 77.415 4.600 77.575 4.700 ;
  LAYER VI1 ;
  RECT 77.445 4.600 77.545 4.700 ;
  LAYER VI2 ;
  RECT 77.445 4.600 77.545 4.700 ;
  LAYER VI3 ;
  RECT 77.445 4.600 77.545 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[34]
PIN DO[34]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 78.815 4.600 78.975 4.700 ;
  LAYER ME2 ;
  RECT 78.815 4.600 78.975 4.700 ;
  LAYER ME1 ;
  RECT 78.815 4.600 78.975 4.700 ;
  LAYER VI1 ;
  RECT 78.845 4.600 78.945 4.700 ;
  LAYER VI2 ;
  RECT 78.845 4.600 78.945 4.700 ;
  LAYER VI3 ;
  RECT 78.845 4.600 78.945 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[34]
PIN DI[33]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 75.315 4.600 75.475 4.700 ;
  LAYER ME2 ;
  RECT 75.315 4.600 75.475 4.700 ;
  LAYER ME1 ;
  RECT 75.315 4.600 75.475 4.700 ;
  LAYER VI1 ;
  RECT 75.345 4.600 75.445 4.700 ;
  LAYER VI2 ;
  RECT 75.345 4.600 75.445 4.700 ;
  LAYER VI3 ;
  RECT 75.345 4.600 75.445 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[33]
PIN DO[33]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 76.715 4.600 76.875 4.700 ;
  LAYER ME2 ;
  RECT 76.715 4.600 76.875 4.700 ;
  LAYER ME1 ;
  RECT 76.715 4.600 76.875 4.700 ;
  LAYER VI1 ;
  RECT 76.745 4.600 76.845 4.700 ;
  LAYER VI2 ;
  RECT 76.745 4.600 76.845 4.700 ;
  LAYER VI3 ;
  RECT 76.745 4.600 76.845 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[33]
PIN DI[32]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 73.215 4.600 73.375 4.700 ;
  LAYER ME2 ;
  RECT 73.215 4.600 73.375 4.700 ;
  LAYER ME1 ;
  RECT 73.215 4.600 73.375 4.700 ;
  LAYER VI1 ;
  RECT 73.245 4.600 73.345 4.700 ;
  LAYER VI2 ;
  RECT 73.245 4.600 73.345 4.700 ;
  LAYER VI3 ;
  RECT 73.245 4.600 73.345 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.088 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.464 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       25.188 LAYER ME2 ;
 ANTENNAMAXAREACAR                       27.726 LAYER ME3 ;
END DI[32]
PIN DO[32]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 74.615 4.600 74.775 4.700 ;
  LAYER ME2 ;
  RECT 74.615 4.600 74.775 4.700 ;
  LAYER ME1 ;
  RECT 74.615 4.600 74.775 4.700 ;
  LAYER VI1 ;
  RECT 74.645 4.600 74.745 4.700 ;
  LAYER VI2 ;
  RECT 74.645 4.600 74.745 4.700 ;
  LAYER VI3 ;
  RECT 74.645 4.600 74.745 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[32]
PIN WEB[1]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 73.485 4.600 73.645 4.700 ;
  LAYER ME2 ;
  RECT 73.485 4.600 73.645 4.700 ;
  LAYER ME1 ;
  RECT 73.485 4.600 73.645 4.700 ;
  LAYER VI1 ;
  RECT 73.515 4.600 73.615 4.700 ;
  LAYER VI2 ;
  RECT 73.515 4.600 73.615 4.700 ;
  LAYER VI3 ;
  RECT 73.515 4.600 73.615 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.093 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.124 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.588 LAYER ME2 ;
 ANTENNAGATEAREA                          0.588 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                        0.618 LAYER ME2 ;
 ANTENNAMAXAREACAR                        0.708 LAYER ME3 ;
END WEB[1]
PIN DI[31]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 71.115 4.600 71.275 4.700 ;
  LAYER ME2 ;
  RECT 71.115 4.600 71.275 4.700 ;
  LAYER ME1 ;
  RECT 71.115 4.600 71.275 4.700 ;
  LAYER VI1 ;
  RECT 71.145 4.600 71.245 4.700 ;
  LAYER VI2 ;
  RECT 71.145 4.600 71.245 4.700 ;
  LAYER VI3 ;
  RECT 71.145 4.600 71.245 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[31]
PIN DO[31]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 72.515 4.600 72.675 4.700 ;
  LAYER ME2 ;
  RECT 72.515 4.600 72.675 4.700 ;
  LAYER ME1 ;
  RECT 72.515 4.600 72.675 4.700 ;
  LAYER VI1 ;
  RECT 72.545 4.600 72.645 4.700 ;
  LAYER VI2 ;
  RECT 72.545 4.600 72.645 4.700 ;
  LAYER VI3 ;
  RECT 72.545 4.600 72.645 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[31]
PIN DI[30]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 69.015 4.600 69.175 4.700 ;
  LAYER ME2 ;
  RECT 69.015 4.600 69.175 4.700 ;
  LAYER ME1 ;
  RECT 69.015 4.600 69.175 4.700 ;
  LAYER VI1 ;
  RECT 69.045 4.600 69.145 4.700 ;
  LAYER VI2 ;
  RECT 69.045 4.600 69.145 4.700 ;
  LAYER VI3 ;
  RECT 69.045 4.600 69.145 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[30]
PIN DO[30]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 70.415 4.600 70.575 4.700 ;
  LAYER ME2 ;
  RECT 70.415 4.600 70.575 4.700 ;
  LAYER ME1 ;
  RECT 70.415 4.600 70.575 4.700 ;
  LAYER VI1 ;
  RECT 70.445 4.600 70.545 4.700 ;
  LAYER VI2 ;
  RECT 70.445 4.600 70.545 4.700 ;
  LAYER VI3 ;
  RECT 70.445 4.600 70.545 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[30]
PIN DI[29]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 66.915 4.600 67.075 4.700 ;
  LAYER ME2 ;
  RECT 66.915 4.600 67.075 4.700 ;
  LAYER ME1 ;
  RECT 66.915 4.600 67.075 4.700 ;
  LAYER VI1 ;
  RECT 66.945 4.600 67.045 4.700 ;
  LAYER VI2 ;
  RECT 66.945 4.600 67.045 4.700 ;
  LAYER VI3 ;
  RECT 66.945 4.600 67.045 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[29]
PIN DO[29]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 68.315 4.600 68.475 4.700 ;
  LAYER ME2 ;
  RECT 68.315 4.600 68.475 4.700 ;
  LAYER ME1 ;
  RECT 68.315 4.600 68.475 4.700 ;
  LAYER VI1 ;
  RECT 68.345 4.600 68.445 4.700 ;
  LAYER VI2 ;
  RECT 68.345 4.600 68.445 4.700 ;
  LAYER VI3 ;
  RECT 68.345 4.600 68.445 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[29]
PIN DI[28]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 64.815 4.600 64.975 4.700 ;
  LAYER ME2 ;
  RECT 64.815 4.600 64.975 4.700 ;
  LAYER ME1 ;
  RECT 64.815 4.600 64.975 4.700 ;
  LAYER VI1 ;
  RECT 64.845 4.600 64.945 4.700 ;
  LAYER VI2 ;
  RECT 64.845 4.600 64.945 4.700 ;
  LAYER VI3 ;
  RECT 64.845 4.600 64.945 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[28]
PIN DO[28]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 66.215 4.600 66.375 4.700 ;
  LAYER ME2 ;
  RECT 66.215 4.600 66.375 4.700 ;
  LAYER ME1 ;
  RECT 66.215 4.600 66.375 4.700 ;
  LAYER VI1 ;
  RECT 66.245 4.600 66.345 4.700 ;
  LAYER VI2 ;
  RECT 66.245 4.600 66.345 4.700 ;
  LAYER VI3 ;
  RECT 66.245 4.600 66.345 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[28]
PIN DI[27]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 62.715 4.600 62.875 4.700 ;
  LAYER ME2 ;
  RECT 62.715 4.600 62.875 4.700 ;
  LAYER ME1 ;
  RECT 62.715 4.600 62.875 4.700 ;
  LAYER VI1 ;
  RECT 62.745 4.600 62.845 4.700 ;
  LAYER VI2 ;
  RECT 62.745 4.600 62.845 4.700 ;
  LAYER VI3 ;
  RECT 62.745 4.600 62.845 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[27]
PIN DO[27]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 64.115 4.600 64.275 4.700 ;
  LAYER ME2 ;
  RECT 64.115 4.600 64.275 4.700 ;
  LAYER ME1 ;
  RECT 64.115 4.600 64.275 4.700 ;
  LAYER VI1 ;
  RECT 64.145 4.600 64.245 4.700 ;
  LAYER VI2 ;
  RECT 64.145 4.600 64.245 4.700 ;
  LAYER VI3 ;
  RECT 64.145 4.600 64.245 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[27]
PIN DI[26]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 60.615 4.600 60.775 4.700 ;
  LAYER ME2 ;
  RECT 60.615 4.600 60.775 4.700 ;
  LAYER ME1 ;
  RECT 60.615 4.600 60.775 4.700 ;
  LAYER VI1 ;
  RECT 60.645 4.600 60.745 4.700 ;
  LAYER VI2 ;
  RECT 60.645 4.600 60.745 4.700 ;
  LAYER VI3 ;
  RECT 60.645 4.600 60.745 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[26]
PIN DO[26]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 62.015 4.600 62.175 4.700 ;
  LAYER ME2 ;
  RECT 62.015 4.600 62.175 4.700 ;
  LAYER ME1 ;
  RECT 62.015 4.600 62.175 4.700 ;
  LAYER VI1 ;
  RECT 62.045 4.600 62.145 4.700 ;
  LAYER VI2 ;
  RECT 62.045 4.600 62.145 4.700 ;
  LAYER VI3 ;
  RECT 62.045 4.600 62.145 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[26]
PIN DI[25]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 58.515 4.600 58.675 4.700 ;
  LAYER ME2 ;
  RECT 58.515 4.600 58.675 4.700 ;
  LAYER ME1 ;
  RECT 58.515 4.600 58.675 4.700 ;
  LAYER VI1 ;
  RECT 58.545 4.600 58.645 4.700 ;
  LAYER VI2 ;
  RECT 58.545 4.600 58.645 4.700 ;
  LAYER VI3 ;
  RECT 58.545 4.600 58.645 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[25]
PIN DO[25]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 59.915 4.600 60.075 4.700 ;
  LAYER ME2 ;
  RECT 59.915 4.600 60.075 4.700 ;
  LAYER ME1 ;
  RECT 59.915 4.600 60.075 4.700 ;
  LAYER VI1 ;
  RECT 59.945 4.600 60.045 4.700 ;
  LAYER VI2 ;
  RECT 59.945 4.600 60.045 4.700 ;
  LAYER VI3 ;
  RECT 59.945 4.600 60.045 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[25]
PIN DI[24]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 56.415 4.600 56.575 4.700 ;
  LAYER ME2 ;
  RECT 56.415 4.600 56.575 4.700 ;
  LAYER ME1 ;
  RECT 56.415 4.600 56.575 4.700 ;
  LAYER VI1 ;
  RECT 56.445 4.600 56.545 4.700 ;
  LAYER VI2 ;
  RECT 56.445 4.600 56.545 4.700 ;
  LAYER VI3 ;
  RECT 56.445 4.600 56.545 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[24]
PIN DO[24]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 57.815 4.600 57.975 4.700 ;
  LAYER ME2 ;
  RECT 57.815 4.600 57.975 4.700 ;
  LAYER ME1 ;
  RECT 57.815 4.600 57.975 4.700 ;
  LAYER VI1 ;
  RECT 57.845 4.600 57.945 4.700 ;
  LAYER VI2 ;
  RECT 57.845 4.600 57.945 4.700 ;
  LAYER VI3 ;
  RECT 57.845 4.600 57.945 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[24]
PIN DI[23]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 54.315 4.600 54.475 4.700 ;
  LAYER ME2 ;
  RECT 54.315 4.600 54.475 4.700 ;
  LAYER ME1 ;
  RECT 54.315 4.600 54.475 4.700 ;
  LAYER VI1 ;
  RECT 54.345 4.600 54.445 4.700 ;
  LAYER VI2 ;
  RECT 54.345 4.600 54.445 4.700 ;
  LAYER VI3 ;
  RECT 54.345 4.600 54.445 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[23]
PIN DO[23]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 55.715 4.600 55.875 4.700 ;
  LAYER ME2 ;
  RECT 55.715 4.600 55.875 4.700 ;
  LAYER ME1 ;
  RECT 55.715 4.600 55.875 4.700 ;
  LAYER VI1 ;
  RECT 55.745 4.600 55.845 4.700 ;
  LAYER VI2 ;
  RECT 55.745 4.600 55.845 4.700 ;
  LAYER VI3 ;
  RECT 55.745 4.600 55.845 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[23]
PIN DI[22]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 52.215 4.600 52.375 4.700 ;
  LAYER ME2 ;
  RECT 52.215 4.600 52.375 4.700 ;
  LAYER ME1 ;
  RECT 52.215 4.600 52.375 4.700 ;
  LAYER VI1 ;
  RECT 52.245 4.600 52.345 4.700 ;
  LAYER VI2 ;
  RECT 52.245 4.600 52.345 4.700 ;
  LAYER VI3 ;
  RECT 52.245 4.600 52.345 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[22]
PIN DO[22]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 53.615 4.600 53.775 4.700 ;
  LAYER ME2 ;
  RECT 53.615 4.600 53.775 4.700 ;
  LAYER ME1 ;
  RECT 53.615 4.600 53.775 4.700 ;
  LAYER VI1 ;
  RECT 53.645 4.600 53.745 4.700 ;
  LAYER VI2 ;
  RECT 53.645 4.600 53.745 4.700 ;
  LAYER VI3 ;
  RECT 53.645 4.600 53.745 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[22]
PIN DI[21]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 50.115 4.600 50.275 4.700 ;
  LAYER ME2 ;
  RECT 50.115 4.600 50.275 4.700 ;
  LAYER ME1 ;
  RECT 50.115 4.600 50.275 4.700 ;
  LAYER VI1 ;
  RECT 50.145 4.600 50.245 4.700 ;
  LAYER VI2 ;
  RECT 50.145 4.600 50.245 4.700 ;
  LAYER VI3 ;
  RECT 50.145 4.600 50.245 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[21]
PIN DO[21]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 51.515 4.600 51.675 4.700 ;
  LAYER ME2 ;
  RECT 51.515 4.600 51.675 4.700 ;
  LAYER ME1 ;
  RECT 51.515 4.600 51.675 4.700 ;
  LAYER VI1 ;
  RECT 51.545 4.600 51.645 4.700 ;
  LAYER VI2 ;
  RECT 51.545 4.600 51.645 4.700 ;
  LAYER VI3 ;
  RECT 51.545 4.600 51.645 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[21]
PIN DI[20]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 48.015 4.600 48.175 4.700 ;
  LAYER ME2 ;
  RECT 48.015 4.600 48.175 4.700 ;
  LAYER ME1 ;
  RECT 48.015 4.600 48.175 4.700 ;
  LAYER VI1 ;
  RECT 48.045 4.600 48.145 4.700 ;
  LAYER VI2 ;
  RECT 48.045 4.600 48.145 4.700 ;
  LAYER VI3 ;
  RECT 48.045 4.600 48.145 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[20]
PIN DO[20]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 49.415 4.600 49.575 4.700 ;
  LAYER ME2 ;
  RECT 49.415 4.600 49.575 4.700 ;
  LAYER ME1 ;
  RECT 49.415 4.600 49.575 4.700 ;
  LAYER VI1 ;
  RECT 49.445 4.600 49.545 4.700 ;
  LAYER VI2 ;
  RECT 49.445 4.600 49.545 4.700 ;
  LAYER VI3 ;
  RECT 49.445 4.600 49.545 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[20]
PIN DI[19]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 45.915 4.600 46.075 4.700 ;
  LAYER ME2 ;
  RECT 45.915 4.600 46.075 4.700 ;
  LAYER ME1 ;
  RECT 45.915 4.600 46.075 4.700 ;
  LAYER VI1 ;
  RECT 45.945 4.600 46.045 4.700 ;
  LAYER VI2 ;
  RECT 45.945 4.600 46.045 4.700 ;
  LAYER VI3 ;
  RECT 45.945 4.600 46.045 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[19]
PIN DO[19]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 47.315 4.600 47.475 4.700 ;
  LAYER ME2 ;
  RECT 47.315 4.600 47.475 4.700 ;
  LAYER ME1 ;
  RECT 47.315 4.600 47.475 4.700 ;
  LAYER VI1 ;
  RECT 47.345 4.600 47.445 4.700 ;
  LAYER VI2 ;
  RECT 47.345 4.600 47.445 4.700 ;
  LAYER VI3 ;
  RECT 47.345 4.600 47.445 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[19]
PIN DI[18]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 43.815 4.600 43.975 4.700 ;
  LAYER ME2 ;
  RECT 43.815 4.600 43.975 4.700 ;
  LAYER ME1 ;
  RECT 43.815 4.600 43.975 4.700 ;
  LAYER VI1 ;
  RECT 43.845 4.600 43.945 4.700 ;
  LAYER VI2 ;
  RECT 43.845 4.600 43.945 4.700 ;
  LAYER VI3 ;
  RECT 43.845 4.600 43.945 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[18]
PIN DO[18]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 45.215 4.600 45.375 4.700 ;
  LAYER ME2 ;
  RECT 45.215 4.600 45.375 4.700 ;
  LAYER ME1 ;
  RECT 45.215 4.600 45.375 4.700 ;
  LAYER VI1 ;
  RECT 45.245 4.600 45.345 4.700 ;
  LAYER VI2 ;
  RECT 45.245 4.600 45.345 4.700 ;
  LAYER VI3 ;
  RECT 45.245 4.600 45.345 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[18]
PIN DI[17]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 41.715 4.600 41.875 4.700 ;
  LAYER ME2 ;
  RECT 41.715 4.600 41.875 4.700 ;
  LAYER ME1 ;
  RECT 41.715 4.600 41.875 4.700 ;
  LAYER VI1 ;
  RECT 41.745 4.600 41.845 4.700 ;
  LAYER VI2 ;
  RECT 41.745 4.600 41.845 4.700 ;
  LAYER VI3 ;
  RECT 41.745 4.600 41.845 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[17]
PIN DO[17]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 43.115 4.600 43.275 4.700 ;
  LAYER ME2 ;
  RECT 43.115 4.600 43.275 4.700 ;
  LAYER ME1 ;
  RECT 43.115 4.600 43.275 4.700 ;
  LAYER VI1 ;
  RECT 43.145 4.600 43.245 4.700 ;
  LAYER VI2 ;
  RECT 43.145 4.600 43.245 4.700 ;
  LAYER VI3 ;
  RECT 43.145 4.600 43.245 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[17]
PIN DI[16]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 39.615 4.600 39.775 4.700 ;
  LAYER ME2 ;
  RECT 39.615 4.600 39.775 4.700 ;
  LAYER ME1 ;
  RECT 39.615 4.600 39.775 4.700 ;
  LAYER VI1 ;
  RECT 39.645 4.600 39.745 4.700 ;
  LAYER VI2 ;
  RECT 39.645 4.600 39.745 4.700 ;
  LAYER VI3 ;
  RECT 39.645 4.600 39.745 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[16]
PIN DO[16]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 41.015 4.600 41.175 4.700 ;
  LAYER ME2 ;
  RECT 41.015 4.600 41.175 4.700 ;
  LAYER ME1 ;
  RECT 41.015 4.600 41.175 4.700 ;
  LAYER VI1 ;
  RECT 41.045 4.600 41.145 4.700 ;
  LAYER VI2 ;
  RECT 41.045 4.600 41.145 4.700 ;
  LAYER VI3 ;
  RECT 41.045 4.600 41.145 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[16]
PIN DI[15]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 37.515 4.600 37.675 4.700 ;
  LAYER ME2 ;
  RECT 37.515 4.600 37.675 4.700 ;
  LAYER ME1 ;
  RECT 37.515 4.600 37.675 4.700 ;
  LAYER VI1 ;
  RECT 37.545 4.600 37.645 4.700 ;
  LAYER VI2 ;
  RECT 37.545 4.600 37.645 4.700 ;
  LAYER VI3 ;
  RECT 37.545 4.600 37.645 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[15]
PIN DO[15]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 38.915 4.600 39.075 4.700 ;
  LAYER ME2 ;
  RECT 38.915 4.600 39.075 4.700 ;
  LAYER ME1 ;
  RECT 38.915 4.600 39.075 4.700 ;
  LAYER VI1 ;
  RECT 38.945 4.600 39.045 4.700 ;
  LAYER VI2 ;
  RECT 38.945 4.600 39.045 4.700 ;
  LAYER VI3 ;
  RECT 38.945 4.600 39.045 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[15]
PIN DI[14]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 35.415 4.600 35.575 4.700 ;
  LAYER ME2 ;
  RECT 35.415 4.600 35.575 4.700 ;
  LAYER ME1 ;
  RECT 35.415 4.600 35.575 4.700 ;
  LAYER VI1 ;
  RECT 35.445 4.600 35.545 4.700 ;
  LAYER VI2 ;
  RECT 35.445 4.600 35.545 4.700 ;
  LAYER VI3 ;
  RECT 35.445 4.600 35.545 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[14]
PIN DO[14]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 36.815 4.600 36.975 4.700 ;
  LAYER ME2 ;
  RECT 36.815 4.600 36.975 4.700 ;
  LAYER ME1 ;
  RECT 36.815 4.600 36.975 4.700 ;
  LAYER VI1 ;
  RECT 36.845 4.600 36.945 4.700 ;
  LAYER VI2 ;
  RECT 36.845 4.600 36.945 4.700 ;
  LAYER VI3 ;
  RECT 36.845 4.600 36.945 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[14]
PIN DI[13]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 33.315 4.600 33.475 4.700 ;
  LAYER ME2 ;
  RECT 33.315 4.600 33.475 4.700 ;
  LAYER ME1 ;
  RECT 33.315 4.600 33.475 4.700 ;
  LAYER VI1 ;
  RECT 33.345 4.600 33.445 4.700 ;
  LAYER VI2 ;
  RECT 33.345 4.600 33.445 4.700 ;
  LAYER VI3 ;
  RECT 33.345 4.600 33.445 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[13]
PIN DO[13]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 34.715 4.600 34.875 4.700 ;
  LAYER ME2 ;
  RECT 34.715 4.600 34.875 4.700 ;
  LAYER ME1 ;
  RECT 34.715 4.600 34.875 4.700 ;
  LAYER VI1 ;
  RECT 34.745 4.600 34.845 4.700 ;
  LAYER VI2 ;
  RECT 34.745 4.600 34.845 4.700 ;
  LAYER VI3 ;
  RECT 34.745 4.600 34.845 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[13]
PIN DI[12]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 31.215 4.600 31.375 4.700 ;
  LAYER ME2 ;
  RECT 31.215 4.600 31.375 4.700 ;
  LAYER ME1 ;
  RECT 31.215 4.600 31.375 4.700 ;
  LAYER VI1 ;
  RECT 31.245 4.600 31.345 4.700 ;
  LAYER VI2 ;
  RECT 31.245 4.600 31.345 4.700 ;
  LAYER VI3 ;
  RECT 31.245 4.600 31.345 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[12]
PIN DO[12]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 32.615 4.600 32.775 4.700 ;
  LAYER ME2 ;
  RECT 32.615 4.600 32.775 4.700 ;
  LAYER ME1 ;
  RECT 32.615 4.600 32.775 4.700 ;
  LAYER VI1 ;
  RECT 32.645 4.600 32.745 4.700 ;
  LAYER VI2 ;
  RECT 32.645 4.600 32.745 4.700 ;
  LAYER VI3 ;
  RECT 32.645 4.600 32.745 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[12]
PIN DI[11]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 29.115 4.600 29.275 4.700 ;
  LAYER ME2 ;
  RECT 29.115 4.600 29.275 4.700 ;
  LAYER ME1 ;
  RECT 29.115 4.600 29.275 4.700 ;
  LAYER VI1 ;
  RECT 29.145 4.600 29.245 4.700 ;
  LAYER VI2 ;
  RECT 29.145 4.600 29.245 4.700 ;
  LAYER VI3 ;
  RECT 29.145 4.600 29.245 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[11]
PIN DO[11]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 30.515 4.600 30.675 4.700 ;
  LAYER ME2 ;
  RECT 30.515 4.600 30.675 4.700 ;
  LAYER ME1 ;
  RECT 30.515 4.600 30.675 4.700 ;
  LAYER VI1 ;
  RECT 30.545 4.600 30.645 4.700 ;
  LAYER VI2 ;
  RECT 30.545 4.600 30.645 4.700 ;
  LAYER VI3 ;
  RECT 30.545 4.600 30.645 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[11]
PIN DI[10]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 27.015 4.600 27.175 4.700 ;
  LAYER ME2 ;
  RECT 27.015 4.600 27.175 4.700 ;
  LAYER ME1 ;
  RECT 27.015 4.600 27.175 4.700 ;
  LAYER VI1 ;
  RECT 27.045 4.600 27.145 4.700 ;
  LAYER VI2 ;
  RECT 27.045 4.600 27.145 4.700 ;
  LAYER VI3 ;
  RECT 27.045 4.600 27.145 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[10]
PIN DO[10]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 28.415 4.600 28.575 4.700 ;
  LAYER ME2 ;
  RECT 28.415 4.600 28.575 4.700 ;
  LAYER ME1 ;
  RECT 28.415 4.600 28.575 4.700 ;
  LAYER VI1 ;
  RECT 28.445 4.600 28.545 4.700 ;
  LAYER VI2 ;
  RECT 28.445 4.600 28.545 4.700 ;
  LAYER VI3 ;
  RECT 28.445 4.600 28.545 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[10]
PIN DI[9]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 24.915 4.600 25.075 4.700 ;
  LAYER ME2 ;
  RECT 24.915 4.600 25.075 4.700 ;
  LAYER ME1 ;
  RECT 24.915 4.600 25.075 4.700 ;
  LAYER VI1 ;
  RECT 24.945 4.600 25.045 4.700 ;
  LAYER VI2 ;
  RECT 24.945 4.600 25.045 4.700 ;
  LAYER VI3 ;
  RECT 24.945 4.600 25.045 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[9]
PIN DO[9]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 26.315 4.600 26.475 4.700 ;
  LAYER ME2 ;
  RECT 26.315 4.600 26.475 4.700 ;
  LAYER ME1 ;
  RECT 26.315 4.600 26.475 4.700 ;
  LAYER VI1 ;
  RECT 26.345 4.600 26.445 4.700 ;
  LAYER VI2 ;
  RECT 26.345 4.600 26.445 4.700 ;
  LAYER VI3 ;
  RECT 26.345 4.600 26.445 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[9]
PIN DI[8]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 22.815 4.600 22.975 4.700 ;
  LAYER ME2 ;
  RECT 22.815 4.600 22.975 4.700 ;
  LAYER ME1 ;
  RECT 22.815 4.600 22.975 4.700 ;
  LAYER VI1 ;
  RECT 22.845 4.600 22.945 4.700 ;
  LAYER VI2 ;
  RECT 22.845 4.600 22.945 4.700 ;
  LAYER VI3 ;
  RECT 22.845 4.600 22.945 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[8]
PIN DO[8]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 24.215 4.600 24.375 4.700 ;
  LAYER ME2 ;
  RECT 24.215 4.600 24.375 4.700 ;
  LAYER ME1 ;
  RECT 24.215 4.600 24.375 4.700 ;
  LAYER VI1 ;
  RECT 24.245 4.600 24.345 4.700 ;
  LAYER VI2 ;
  RECT 24.245 4.600 24.345 4.700 ;
  LAYER VI3 ;
  RECT 24.245 4.600 24.345 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[8]
PIN DI[7]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 20.715 4.600 20.875 4.700 ;
  LAYER ME2 ;
  RECT 20.715 4.600 20.875 4.700 ;
  LAYER ME1 ;
  RECT 20.715 4.600 20.875 4.700 ;
  LAYER VI1 ;
  RECT 20.745 4.600 20.845 4.700 ;
  LAYER VI2 ;
  RECT 20.745 4.600 20.845 4.700 ;
  LAYER VI3 ;
  RECT 20.745 4.600 20.845 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[7]
PIN DO[7]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 22.115 4.600 22.275 4.700 ;
  LAYER ME2 ;
  RECT 22.115 4.600 22.275 4.700 ;
  LAYER ME1 ;
  RECT 22.115 4.600 22.275 4.700 ;
  LAYER VI1 ;
  RECT 22.145 4.600 22.245 4.700 ;
  LAYER VI2 ;
  RECT 22.145 4.600 22.245 4.700 ;
  LAYER VI3 ;
  RECT 22.145 4.600 22.245 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[7]
PIN DI[6]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 18.615 4.600 18.775 4.700 ;
  LAYER ME2 ;
  RECT 18.615 4.600 18.775 4.700 ;
  LAYER ME1 ;
  RECT 18.615 4.600 18.775 4.700 ;
  LAYER VI1 ;
  RECT 18.645 4.600 18.745 4.700 ;
  LAYER VI2 ;
  RECT 18.645 4.600 18.745 4.700 ;
  LAYER VI3 ;
  RECT 18.645 4.600 18.745 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[6]
PIN DO[6]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 20.015 4.600 20.175 4.700 ;
  LAYER ME2 ;
  RECT 20.015 4.600 20.175 4.700 ;
  LAYER ME1 ;
  RECT 20.015 4.600 20.175 4.700 ;
  LAYER VI1 ;
  RECT 20.045 4.600 20.145 4.700 ;
  LAYER VI2 ;
  RECT 20.045 4.600 20.145 4.700 ;
  LAYER VI3 ;
  RECT 20.045 4.600 20.145 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[6]
PIN DI[5]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 16.515 4.600 16.675 4.700 ;
  LAYER ME2 ;
  RECT 16.515 4.600 16.675 4.700 ;
  LAYER ME1 ;
  RECT 16.515 4.600 16.675 4.700 ;
  LAYER VI1 ;
  RECT 16.545 4.600 16.645 4.700 ;
  LAYER VI2 ;
  RECT 16.545 4.600 16.645 4.700 ;
  LAYER VI3 ;
  RECT 16.545 4.600 16.645 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[5]
PIN DO[5]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 17.915 4.600 18.075 4.700 ;
  LAYER ME2 ;
  RECT 17.915 4.600 18.075 4.700 ;
  LAYER ME1 ;
  RECT 17.915 4.600 18.075 4.700 ;
  LAYER VI1 ;
  RECT 17.945 4.600 18.045 4.700 ;
  LAYER VI2 ;
  RECT 17.945 4.600 18.045 4.700 ;
  LAYER VI3 ;
  RECT 17.945 4.600 18.045 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[5]
PIN DI[4]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 14.415 4.600 14.575 4.700 ;
  LAYER ME2 ;
  RECT 14.415 4.600 14.575 4.700 ;
  LAYER ME1 ;
  RECT 14.415 4.600 14.575 4.700 ;
  LAYER VI1 ;
  RECT 14.445 4.600 14.545 4.700 ;
  LAYER VI2 ;
  RECT 14.445 4.600 14.545 4.700 ;
  LAYER VI3 ;
  RECT 14.445 4.600 14.545 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[4]
PIN DO[4]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 15.815 4.600 15.975 4.700 ;
  LAYER ME2 ;
  RECT 15.815 4.600 15.975 4.700 ;
  LAYER ME1 ;
  RECT 15.815 4.600 15.975 4.700 ;
  LAYER VI1 ;
  RECT 15.845 4.600 15.945 4.700 ;
  LAYER VI2 ;
  RECT 15.845 4.600 15.945 4.700 ;
  LAYER VI3 ;
  RECT 15.845 4.600 15.945 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[4]
PIN DI[3]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 12.315 4.600 12.475 4.700 ;
  LAYER ME2 ;
  RECT 12.315 4.600 12.475 4.700 ;
  LAYER ME1 ;
  RECT 12.315 4.600 12.475 4.700 ;
  LAYER VI1 ;
  RECT 12.345 4.600 12.445 4.700 ;
  LAYER VI2 ;
  RECT 12.345 4.600 12.445 4.700 ;
  LAYER VI3 ;
  RECT 12.345 4.600 12.445 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[3]
PIN DO[3]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 13.715 4.600 13.875 4.700 ;
  LAYER ME2 ;
  RECT 13.715 4.600 13.875 4.700 ;
  LAYER ME1 ;
  RECT 13.715 4.600 13.875 4.700 ;
  LAYER VI1 ;
  RECT 13.745 4.600 13.845 4.700 ;
  LAYER VI2 ;
  RECT 13.745 4.600 13.845 4.700 ;
  LAYER VI3 ;
  RECT 13.745 4.600 13.845 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[3]
PIN DI[2]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 10.215 4.600 10.375 4.700 ;
  LAYER ME2 ;
  RECT 10.215 4.600 10.375 4.700 ;
  LAYER ME1 ;
  RECT 10.215 4.600 10.375 4.700 ;
  LAYER VI1 ;
  RECT 10.245 4.600 10.345 4.700 ;
  LAYER VI2 ;
  RECT 10.245 4.600 10.345 4.700 ;
  LAYER VI3 ;
  RECT 10.245 4.600 10.345 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[2]
PIN DO[2]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 11.615 4.600 11.775 4.700 ;
  LAYER ME2 ;
  RECT 11.615 4.600 11.775 4.700 ;
  LAYER ME1 ;
  RECT 11.615 4.600 11.775 4.700 ;
  LAYER VI1 ;
  RECT 11.645 4.600 11.745 4.700 ;
  LAYER VI2 ;
  RECT 11.645 4.600 11.745 4.700 ;
  LAYER VI3 ;
  RECT 11.645 4.600 11.745 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[2]
PIN DI[1]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 8.115 4.600 8.275 4.700 ;
  LAYER ME2 ;
  RECT 8.115 4.600 8.275 4.700 ;
  LAYER ME1 ;
  RECT 8.115 4.600 8.275 4.700 ;
  LAYER VI1 ;
  RECT 8.145 4.600 8.245 4.700 ;
  LAYER VI2 ;
  RECT 8.145 4.600 8.245 4.700 ;
  LAYER VI3 ;
  RECT 8.145 4.600 8.245 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[1]
PIN DO[1]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 9.515 4.600 9.675 4.700 ;
  LAYER ME2 ;
  RECT 9.515 4.600 9.675 4.700 ;
  LAYER ME1 ;
  RECT 9.515 4.600 9.675 4.700 ;
  LAYER VI1 ;
  RECT 9.545 4.600 9.645 4.700 ;
  LAYER VI2 ;
  RECT 9.545 4.600 9.645 4.700 ;
  LAYER VI3 ;
  RECT 9.545 4.600 9.645 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[1]
PIN DI[0]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 6.015 4.600 6.175 4.700 ;
  LAYER ME2 ;
  RECT 6.015 4.600 6.175 4.700 ;
  LAYER ME1 ;
  RECT 6.015 4.600 6.175 4.700 ;
  LAYER VI1 ;
  RECT 6.045 4.600 6.145 4.700 ;
  LAYER VI2 ;
  RECT 6.045 4.600 6.145 4.700 ;
  LAYER VI3 ;
  RECT 6.045 4.600 6.145 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.088 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.464 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       25.188 LAYER ME2 ;
 ANTENNAMAXAREACAR                       27.726 LAYER ME3 ;
END DI[0]
PIN DO[0]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 7.415 4.600 7.575 4.700 ;
  LAYER ME2 ;
  RECT 7.415 4.600 7.575 4.700 ;
  LAYER ME1 ;
  RECT 7.415 4.600 7.575 4.700 ;
  LAYER VI1 ;
  RECT 7.445 4.600 7.545 4.700 ;
  LAYER VI2 ;
  RECT 7.445 4.600 7.545 4.700 ;
  LAYER VI3 ;
  RECT 7.445 4.600 7.545 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[0]
PIN WEB[0]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 6.285 4.600 6.445 4.700 ;
  LAYER ME2 ;
  RECT 6.285 4.600 6.445 4.700 ;
  LAYER ME1 ;
  RECT 6.285 4.600 6.445 4.700 ;
  LAYER VI1 ;
  RECT 6.315 4.600 6.415 4.700 ;
  LAYER VI2 ;
  RECT 6.315 4.600 6.415 4.700 ;
  LAYER VI3 ;
  RECT 6.315 4.600 6.415 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.093 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.124 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.588 LAYER ME2 ;
 ANTENNAGATEAREA                          0.588 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                        0.618 LAYER ME2 ;
 ANTENNAMAXAREACAR                        0.708 LAYER ME3 ;
END WEB[0]
PIN A[8]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 141.235 4.600 141.395 4.750 ;
  LAYER ME2 ;
  RECT 141.235 4.600 141.395 4.750 ;
  LAYER ME1 ;
  RECT 141.235 4.600 141.395 4.750 ;
  LAYER VI1 ;
  RECT 141.265 4.600 141.365 4.700 ;
  LAYER VI2 ;
  RECT 141.265 4.600 141.365 4.700 ;
  LAYER VI3 ;
  RECT 141.265 4.600 141.365 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.029 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  1.277 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.029 LAYER ME3 ;
 ANTENNAGATEAREA                          0.138 LAYER ME2 ;
 ANTENNAGATEAREA                          0.138 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                        9.783 LAYER ME2 ;
 ANTENNAMAXAREACAR                       10.166 LAYER ME3 ;
END A[8]
PIN A[7]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 142.320 4.600 142.480 4.750 ;
  LAYER ME2 ;
  RECT 142.320 4.600 142.480 4.750 ;
  LAYER ME1 ;
  RECT 142.320 4.600 142.480 4.750 ;
  LAYER VI1 ;
  RECT 142.350 4.600 142.450 4.700 ;
  LAYER VI2 ;
  RECT 142.350 4.600 142.450 4.700 ;
  LAYER VI3 ;
  RECT 142.350 4.600 142.450 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.029 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  1.296 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.029 LAYER ME3 ;
 ANTENNAGATEAREA                          0.138 LAYER ME2 ;
 ANTENNAGATEAREA                          0.138 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                        9.917 LAYER ME2 ;
 ANTENNAMAXAREACAR                       10.300 LAYER ME3 ;
END A[7]
PIN A[6]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 143.515 4.600 143.675 4.750 ;
  LAYER ME2 ;
  RECT 143.515 4.600 143.675 4.750 ;
  LAYER ME1 ;
  RECT 143.515 4.600 143.675 4.750 ;
  LAYER VI1 ;
  RECT 143.545 4.600 143.645 4.700 ;
  LAYER VI2 ;
  RECT 143.545 4.600 143.645 4.700 ;
  LAYER VI3 ;
  RECT 143.545 4.600 143.645 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.029 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  1.277 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.029 LAYER ME3 ;
 ANTENNAGATEAREA                          0.138 LAYER ME2 ;
 ANTENNAGATEAREA                          0.138 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                        9.783 LAYER ME2 ;
 ANTENNAMAXAREACAR                       10.166 LAYER ME3 ;
END A[6]
PIN A[5]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 144.600 4.600 144.760 4.750 ;
  LAYER ME2 ;
  RECT 144.600 4.600 144.760 4.750 ;
  LAYER ME1 ;
  RECT 144.600 4.600 144.760 4.750 ;
  LAYER VI1 ;
  RECT 144.630 4.600 144.730 4.700 ;
  LAYER VI2 ;
  RECT 144.630 4.600 144.730 4.700 ;
  LAYER VI3 ;
  RECT 144.630 4.600 144.730 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.029 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  1.296 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.029 LAYER ME3 ;
 ANTENNAGATEAREA                          0.138 LAYER ME2 ;
 ANTENNAGATEAREA                          0.138 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                        9.917 LAYER ME2 ;
 ANTENNAMAXAREACAR                       10.300 LAYER ME3 ;
END A[5]
PIN A[4]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 145.795 4.600 145.955 4.750 ;
  LAYER ME2 ;
  RECT 145.795 4.600 145.955 4.750 ;
  LAYER ME1 ;
  RECT 145.795 4.600 145.955 4.750 ;
  LAYER VI1 ;
  RECT 145.825 4.600 145.925 4.700 ;
  LAYER VI2 ;
  RECT 145.825 4.600 145.925 4.700 ;
  LAYER VI3 ;
  RECT 145.825 4.600 145.925 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.029 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  1.277 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.029 LAYER ME3 ;
 ANTENNAGATEAREA                          0.138 LAYER ME2 ;
 ANTENNAGATEAREA                          0.138 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                        9.783 LAYER ME2 ;
 ANTENNAMAXAREACAR                       10.166 LAYER ME3 ;
END A[4]
PIN A[3]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 146.880 4.600 147.040 4.750 ;
  LAYER ME2 ;
  RECT 146.880 4.600 147.040 4.750 ;
  LAYER ME1 ;
  RECT 146.880 4.600 147.040 4.750 ;
  LAYER VI1 ;
  RECT 146.910 4.600 147.010 4.700 ;
  LAYER VI2 ;
  RECT 146.910 4.600 147.010 4.700 ;
  LAYER VI3 ;
  RECT 146.910 4.600 147.010 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.029 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  1.296 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.029 LAYER ME3 ;
 ANTENNAGATEAREA                          0.138 LAYER ME2 ;
 ANTENNAGATEAREA                          0.138 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                        9.917 LAYER ME2 ;
 ANTENNAMAXAREACAR                       10.300 LAYER ME3 ;
END A[3]
PIN A[2]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 147.780 4.600 147.940 4.770 ;
  LAYER ME2 ;
  RECT 147.780 4.600 147.940 4.770 ;
  LAYER ME1 ;
  RECT 147.780 4.600 147.940 4.770 ;
  LAYER VI1 ;
  RECT 147.810 4.600 147.910 4.700 ;
  LAYER VI2 ;
  RECT 147.810 4.600 147.910 4.700 ;
  LAYER VI3 ;
  RECT 147.810 4.600 147.910 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.026 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  1.241 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.026 LAYER ME3 ;
 ANTENNAGATEAREA                          0.138 LAYER ME2 ;
 ANTENNAGATEAREA                          0.138 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                        9.548 LAYER ME2 ;
 ANTENNAMAXAREACAR                        9.930 LAYER ME3 ;
END A[2]
PIN A[1]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 148.645 4.600 148.805 4.770 ;
  LAYER ME2 ;
  RECT 148.645 4.600 148.805 4.770 ;
  LAYER ME1 ;
  RECT 148.645 4.600 148.805 4.770 ;
  LAYER VI1 ;
  RECT 148.675 4.600 148.775 4.700 ;
  LAYER VI2 ;
  RECT 148.675 4.600 148.775 4.700 ;
  LAYER VI3 ;
  RECT 148.675 4.600 148.775 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.026 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  1.307 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.026 LAYER ME3 ;
 ANTENNAGATEAREA                          0.138 LAYER ME2 ;
 ANTENNAGATEAREA                          0.138 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       10.025 LAYER ME2 ;
 ANTENNAMAXAREACAR                       10.407 LAYER ME3 ;
END A[1]
PIN A[0]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 151.085 4.600 151.245 4.750 ;
  LAYER ME2 ;
  RECT 151.085 4.600 151.245 4.750 ;
  LAYER ME1 ;
  RECT 151.085 4.600 151.245 4.750 ;
  LAYER VI1 ;
  RECT 151.115 4.600 151.215 4.700 ;
  LAYER VI2 ;
  RECT 151.115 4.600 151.215 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.029 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  1.231 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.029 LAYER ME3 ;
 ANTENNAGATEAREA                          0.138 LAYER ME2 ;
 ANTENNAGATEAREA                          0.138 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                        9.457 LAYER ME2 ;
 ANTENNAMAXAREACAR                        9.839 LAYER ME3 ;
END A[0]
PIN DVSE
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 156.715 4.600 156.875 4.750 ;
  LAYER ME2 ;
  RECT 156.715 4.600 156.875 4.750 ;
  LAYER ME1 ;
  RECT 156.715 4.600 156.875 4.750 ;
  LAYER VI1 ;
  RECT 156.745 4.600 156.845 4.700 ;
  LAYER VI2 ;
  RECT 156.745 4.600 156.845 4.700 ;
  LAYER VI3 ;
  RECT 156.745 4.600 156.845 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.029 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  2.301 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.273 LAYER ME3 ;
 ANTENNAGATEAREA                          0.090 LAYER ME2 ;
 ANTENNAGATEAREA                          0.162 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       26.321 LAYER ME2 ;
 ANTENNAMAXAREACAR                       29.619 LAYER ME3 ;
END DVSE
PIN DVS[3]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 156.175 4.600 156.335 4.750 ;
  LAYER ME2 ;
  RECT 156.175 4.600 156.335 4.750 ;
  LAYER ME1 ;
  RECT 156.175 4.600 156.335 4.750 ;
  LAYER VI1 ;
  RECT 156.205 4.600 156.305 4.700 ;
  LAYER VI2 ;
  RECT 156.205 4.600 156.305 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.029 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  1.802 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.029 LAYER ME3 ;
 ANTENNAGATEAREA                          0.018 LAYER ME2 ;
 ANTENNAGATEAREA                          0.018 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                      105.822 LAYER ME2 ;
 ANTENNAMAXAREACAR                      108.756 LAYER ME3 ;
END DVS[3]
PIN DVS[2]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 156.445 4.600 156.605 4.750 ;
  LAYER ME2 ;
  RECT 156.445 4.600 156.605 4.750 ;
  LAYER ME1 ;
  RECT 156.445 4.600 156.605 4.750 ;
  LAYER VI1 ;
  RECT 156.475 4.600 156.575 4.700 ;
  LAYER VI2 ;
  RECT 156.475 4.600 156.575 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.029 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  1.795 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.029 LAYER ME3 ;
 ANTENNAGATEAREA                          0.018 LAYER ME2 ;
 ANTENNAGATEAREA                          0.018 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                      103.844 LAYER ME2 ;
 ANTENNAMAXAREACAR                      106.778 LAYER ME3 ;
END DVS[2]
PIN DVS[1]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 157.165 4.600 157.325 4.750 ;
  LAYER ME2 ;
  RECT 157.165 4.600 157.325 4.750 ;
  LAYER ME1 ;
  RECT 157.165 4.600 157.325 4.750 ;
  LAYER VI1 ;
  RECT 157.195 4.600 157.295 4.700 ;
  LAYER VI2 ;
  RECT 157.195 4.600 157.295 4.700 ;
  LAYER VI3 ;
  RECT 157.195 4.600 157.295 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.029 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  1.723 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.029 LAYER ME3 ;
 ANTENNAGATEAREA                          0.018 LAYER ME2 ;
 ANTENNAGATEAREA                          0.018 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                      101.853 LAYER ME2 ;
 ANTENNAMAXAREACAR                      104.786 LAYER ME3 ;
END DVS[1]
PIN DVS[0]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 157.450 4.600 157.610 4.750 ;
  LAYER ME2 ;
  RECT 157.450 4.600 157.610 4.750 ;
  LAYER ME1 ;
  RECT 157.450 4.600 157.610 4.750 ;
  LAYER VI1 ;
  RECT 157.480 4.600 157.580 4.700 ;
  LAYER VI2 ;
  RECT 157.480 4.600 157.580 4.700 ;
  LAYER VI3 ;
  RECT 157.480 4.600 157.580 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.029 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  1.729 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.029 LAYER ME3 ;
 ANTENNAGATEAREA                          0.018 LAYER ME2 ;
 ANTENNAGATEAREA                          0.018 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                      100.700 LAYER ME2 ;
 ANTENNAMAXAREACAR                      103.633 LAYER ME3 ;
END DVS[0]
PIN CK
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 150.705 4.600 150.865 4.750 ;
  LAYER ME2 ;
  RECT 150.705 4.600 150.865 4.750 ;
  LAYER ME1 ;
  RECT 150.705 4.600 150.865 4.750 ;
  LAYER VI1 ;
  RECT 150.735 4.600 150.835 4.700 ;
  LAYER VI2 ;
  RECT 150.735 4.600 150.835 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.029 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  1.121 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  1.181 LAYER ME3 ;
 ANTENNAGATEAREA                          0.048 LAYER ME2 ;
 ANTENNAGATEAREA                          0.256 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       25.648 LAYER ME2 ;
 ANTENNAMAXAREACAR                       88.641 LAYER ME3 ;
END CK
PIN CSB
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 150.015 4.600 150.175 4.750 ;
  LAYER ME2 ;
  RECT 150.015 4.600 150.175 4.750 ;
  LAYER ME1 ;
  RECT 150.015 4.600 150.175 4.750 ;
  LAYER VI1 ;
  RECT 150.045 4.600 150.145 4.700 ;
  LAYER VI2 ;
  RECT 150.045 4.600 150.145 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.029 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  1.000 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  1.284 LAYER ME3 ;
 ANTENNAGATEAREA                          0.048 LAYER ME2 ;
 ANTENNAGATEAREA                          0.750 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.308 LAYER ME2 ;
 ANTENNAMAXAREACAR                       49.567 LAYER ME3 ;
END CSB
PIN DI[127]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 290.540 4.600 290.700 4.700 ;
  LAYER ME2 ;
  RECT 290.540 4.600 290.700 4.700 ;
  LAYER ME1 ;
  RECT 290.540 4.600 290.700 4.700 ;
  LAYER VI1 ;
  RECT 290.570 4.600 290.670 4.700 ;
  LAYER VI2 ;
  RECT 290.570 4.600 290.670 4.700 ;
  LAYER VI3 ;
  RECT 290.570 4.600 290.670 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[127]
PIN DO[127]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 291.940 4.600 292.100 4.700 ;
  LAYER ME2 ;
  RECT 291.940 4.600 292.100 4.700 ;
  LAYER ME1 ;
  RECT 291.940 4.600 292.100 4.700 ;
  LAYER VI1 ;
  RECT 291.970 4.600 292.070 4.700 ;
  LAYER VI2 ;
  RECT 291.970 4.600 292.070 4.700 ;
  LAYER VI3 ;
  RECT 291.970 4.600 292.070 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[127]
PIN DI[126]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 288.440 4.600 288.600 4.700 ;
  LAYER ME2 ;
  RECT 288.440 4.600 288.600 4.700 ;
  LAYER ME1 ;
  RECT 288.440 4.600 288.600 4.700 ;
  LAYER VI1 ;
  RECT 288.470 4.600 288.570 4.700 ;
  LAYER VI2 ;
  RECT 288.470 4.600 288.570 4.700 ;
  LAYER VI3 ;
  RECT 288.470 4.600 288.570 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[126]
PIN DO[126]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 289.840 4.600 290.000 4.700 ;
  LAYER ME2 ;
  RECT 289.840 4.600 290.000 4.700 ;
  LAYER ME1 ;
  RECT 289.840 4.600 290.000 4.700 ;
  LAYER VI1 ;
  RECT 289.870 4.600 289.970 4.700 ;
  LAYER VI2 ;
  RECT 289.870 4.600 289.970 4.700 ;
  LAYER VI3 ;
  RECT 289.870 4.600 289.970 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[126]
PIN DI[125]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 286.340 4.600 286.500 4.700 ;
  LAYER ME2 ;
  RECT 286.340 4.600 286.500 4.700 ;
  LAYER ME1 ;
  RECT 286.340 4.600 286.500 4.700 ;
  LAYER VI1 ;
  RECT 286.370 4.600 286.470 4.700 ;
  LAYER VI2 ;
  RECT 286.370 4.600 286.470 4.700 ;
  LAYER VI3 ;
  RECT 286.370 4.600 286.470 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[125]
PIN DO[125]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 287.740 4.600 287.900 4.700 ;
  LAYER ME2 ;
  RECT 287.740 4.600 287.900 4.700 ;
  LAYER ME1 ;
  RECT 287.740 4.600 287.900 4.700 ;
  LAYER VI1 ;
  RECT 287.770 4.600 287.870 4.700 ;
  LAYER VI2 ;
  RECT 287.770 4.600 287.870 4.700 ;
  LAYER VI3 ;
  RECT 287.770 4.600 287.870 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[125]
PIN DI[124]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 284.240 4.600 284.400 4.700 ;
  LAYER ME2 ;
  RECT 284.240 4.600 284.400 4.700 ;
  LAYER ME1 ;
  RECT 284.240 4.600 284.400 4.700 ;
  LAYER VI1 ;
  RECT 284.270 4.600 284.370 4.700 ;
  LAYER VI2 ;
  RECT 284.270 4.600 284.370 4.700 ;
  LAYER VI3 ;
  RECT 284.270 4.600 284.370 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[124]
PIN DO[124]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 285.640 4.600 285.800 4.700 ;
  LAYER ME2 ;
  RECT 285.640 4.600 285.800 4.700 ;
  LAYER ME1 ;
  RECT 285.640 4.600 285.800 4.700 ;
  LAYER VI1 ;
  RECT 285.670 4.600 285.770 4.700 ;
  LAYER VI2 ;
  RECT 285.670 4.600 285.770 4.700 ;
  LAYER VI3 ;
  RECT 285.670 4.600 285.770 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[124]
PIN DI[123]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 282.140 4.600 282.300 4.700 ;
  LAYER ME2 ;
  RECT 282.140 4.600 282.300 4.700 ;
  LAYER ME1 ;
  RECT 282.140 4.600 282.300 4.700 ;
  LAYER VI1 ;
  RECT 282.170 4.600 282.270 4.700 ;
  LAYER VI2 ;
  RECT 282.170 4.600 282.270 4.700 ;
  LAYER VI3 ;
  RECT 282.170 4.600 282.270 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[123]
PIN DO[123]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 283.540 4.600 283.700 4.700 ;
  LAYER ME2 ;
  RECT 283.540 4.600 283.700 4.700 ;
  LAYER ME1 ;
  RECT 283.540 4.600 283.700 4.700 ;
  LAYER VI1 ;
  RECT 283.570 4.600 283.670 4.700 ;
  LAYER VI2 ;
  RECT 283.570 4.600 283.670 4.700 ;
  LAYER VI3 ;
  RECT 283.570 4.600 283.670 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[123]
PIN DI[122]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 280.040 4.600 280.200 4.700 ;
  LAYER ME2 ;
  RECT 280.040 4.600 280.200 4.700 ;
  LAYER ME1 ;
  RECT 280.040 4.600 280.200 4.700 ;
  LAYER VI1 ;
  RECT 280.070 4.600 280.170 4.700 ;
  LAYER VI2 ;
  RECT 280.070 4.600 280.170 4.700 ;
  LAYER VI3 ;
  RECT 280.070 4.600 280.170 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[122]
PIN DO[122]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 281.440 4.600 281.600 4.700 ;
  LAYER ME2 ;
  RECT 281.440 4.600 281.600 4.700 ;
  LAYER ME1 ;
  RECT 281.440 4.600 281.600 4.700 ;
  LAYER VI1 ;
  RECT 281.470 4.600 281.570 4.700 ;
  LAYER VI2 ;
  RECT 281.470 4.600 281.570 4.700 ;
  LAYER VI3 ;
  RECT 281.470 4.600 281.570 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[122]
PIN DI[121]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 277.940 4.600 278.100 4.700 ;
  LAYER ME2 ;
  RECT 277.940 4.600 278.100 4.700 ;
  LAYER ME1 ;
  RECT 277.940 4.600 278.100 4.700 ;
  LAYER VI1 ;
  RECT 277.970 4.600 278.070 4.700 ;
  LAYER VI2 ;
  RECT 277.970 4.600 278.070 4.700 ;
  LAYER VI3 ;
  RECT 277.970 4.600 278.070 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[121]
PIN DO[121]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 279.340 4.600 279.500 4.700 ;
  LAYER ME2 ;
  RECT 279.340 4.600 279.500 4.700 ;
  LAYER ME1 ;
  RECT 279.340 4.600 279.500 4.700 ;
  LAYER VI1 ;
  RECT 279.370 4.600 279.470 4.700 ;
  LAYER VI2 ;
  RECT 279.370 4.600 279.470 4.700 ;
  LAYER VI3 ;
  RECT 279.370 4.600 279.470 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[121]
PIN DI[120]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 275.840 4.600 276.000 4.700 ;
  LAYER ME2 ;
  RECT 275.840 4.600 276.000 4.700 ;
  LAYER ME1 ;
  RECT 275.840 4.600 276.000 4.700 ;
  LAYER VI1 ;
  RECT 275.870 4.600 275.970 4.700 ;
  LAYER VI2 ;
  RECT 275.870 4.600 275.970 4.700 ;
  LAYER VI3 ;
  RECT 275.870 4.600 275.970 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[120]
PIN DO[120]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 277.240 4.600 277.400 4.700 ;
  LAYER ME2 ;
  RECT 277.240 4.600 277.400 4.700 ;
  LAYER ME1 ;
  RECT 277.240 4.600 277.400 4.700 ;
  LAYER VI1 ;
  RECT 277.270 4.600 277.370 4.700 ;
  LAYER VI2 ;
  RECT 277.270 4.600 277.370 4.700 ;
  LAYER VI3 ;
  RECT 277.270 4.600 277.370 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[120]
PIN DI[119]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 273.740 4.600 273.900 4.700 ;
  LAYER ME2 ;
  RECT 273.740 4.600 273.900 4.700 ;
  LAYER ME1 ;
  RECT 273.740 4.600 273.900 4.700 ;
  LAYER VI1 ;
  RECT 273.770 4.600 273.870 4.700 ;
  LAYER VI2 ;
  RECT 273.770 4.600 273.870 4.700 ;
  LAYER VI3 ;
  RECT 273.770 4.600 273.870 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[119]
PIN DO[119]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 275.140 4.600 275.300 4.700 ;
  LAYER ME2 ;
  RECT 275.140 4.600 275.300 4.700 ;
  LAYER ME1 ;
  RECT 275.140 4.600 275.300 4.700 ;
  LAYER VI1 ;
  RECT 275.170 4.600 275.270 4.700 ;
  LAYER VI2 ;
  RECT 275.170 4.600 275.270 4.700 ;
  LAYER VI3 ;
  RECT 275.170 4.600 275.270 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[119]
PIN DI[118]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 271.640 4.600 271.800 4.700 ;
  LAYER ME2 ;
  RECT 271.640 4.600 271.800 4.700 ;
  LAYER ME1 ;
  RECT 271.640 4.600 271.800 4.700 ;
  LAYER VI1 ;
  RECT 271.670 4.600 271.770 4.700 ;
  LAYER VI2 ;
  RECT 271.670 4.600 271.770 4.700 ;
  LAYER VI3 ;
  RECT 271.670 4.600 271.770 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[118]
PIN DO[118]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 273.040 4.600 273.200 4.700 ;
  LAYER ME2 ;
  RECT 273.040 4.600 273.200 4.700 ;
  LAYER ME1 ;
  RECT 273.040 4.600 273.200 4.700 ;
  LAYER VI1 ;
  RECT 273.070 4.600 273.170 4.700 ;
  LAYER VI2 ;
  RECT 273.070 4.600 273.170 4.700 ;
  LAYER VI3 ;
  RECT 273.070 4.600 273.170 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[118]
PIN DI[117]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 269.540 4.600 269.700 4.700 ;
  LAYER ME2 ;
  RECT 269.540 4.600 269.700 4.700 ;
  LAYER ME1 ;
  RECT 269.540 4.600 269.700 4.700 ;
  LAYER VI1 ;
  RECT 269.570 4.600 269.670 4.700 ;
  LAYER VI2 ;
  RECT 269.570 4.600 269.670 4.700 ;
  LAYER VI3 ;
  RECT 269.570 4.600 269.670 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[117]
PIN DO[117]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 270.940 4.600 271.100 4.700 ;
  LAYER ME2 ;
  RECT 270.940 4.600 271.100 4.700 ;
  LAYER ME1 ;
  RECT 270.940 4.600 271.100 4.700 ;
  LAYER VI1 ;
  RECT 270.970 4.600 271.070 4.700 ;
  LAYER VI2 ;
  RECT 270.970 4.600 271.070 4.700 ;
  LAYER VI3 ;
  RECT 270.970 4.600 271.070 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[117]
PIN DI[116]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 267.440 4.600 267.600 4.700 ;
  LAYER ME2 ;
  RECT 267.440 4.600 267.600 4.700 ;
  LAYER ME1 ;
  RECT 267.440 4.600 267.600 4.700 ;
  LAYER VI1 ;
  RECT 267.470 4.600 267.570 4.700 ;
  LAYER VI2 ;
  RECT 267.470 4.600 267.570 4.700 ;
  LAYER VI3 ;
  RECT 267.470 4.600 267.570 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[116]
PIN DO[116]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 268.840 4.600 269.000 4.700 ;
  LAYER ME2 ;
  RECT 268.840 4.600 269.000 4.700 ;
  LAYER ME1 ;
  RECT 268.840 4.600 269.000 4.700 ;
  LAYER VI1 ;
  RECT 268.870 4.600 268.970 4.700 ;
  LAYER VI2 ;
  RECT 268.870 4.600 268.970 4.700 ;
  LAYER VI3 ;
  RECT 268.870 4.600 268.970 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[116]
PIN DI[115]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 265.340 4.600 265.500 4.700 ;
  LAYER ME2 ;
  RECT 265.340 4.600 265.500 4.700 ;
  LAYER ME1 ;
  RECT 265.340 4.600 265.500 4.700 ;
  LAYER VI1 ;
  RECT 265.370 4.600 265.470 4.700 ;
  LAYER VI2 ;
  RECT 265.370 4.600 265.470 4.700 ;
  LAYER VI3 ;
  RECT 265.370 4.600 265.470 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[115]
PIN DO[115]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 266.740 4.600 266.900 4.700 ;
  LAYER ME2 ;
  RECT 266.740 4.600 266.900 4.700 ;
  LAYER ME1 ;
  RECT 266.740 4.600 266.900 4.700 ;
  LAYER VI1 ;
  RECT 266.770 4.600 266.870 4.700 ;
  LAYER VI2 ;
  RECT 266.770 4.600 266.870 4.700 ;
  LAYER VI3 ;
  RECT 266.770 4.600 266.870 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[115]
PIN DI[114]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 263.240 4.600 263.400 4.700 ;
  LAYER ME2 ;
  RECT 263.240 4.600 263.400 4.700 ;
  LAYER ME1 ;
  RECT 263.240 4.600 263.400 4.700 ;
  LAYER VI1 ;
  RECT 263.270 4.600 263.370 4.700 ;
  LAYER VI2 ;
  RECT 263.270 4.600 263.370 4.700 ;
  LAYER VI3 ;
  RECT 263.270 4.600 263.370 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[114]
PIN DO[114]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 264.640 4.600 264.800 4.700 ;
  LAYER ME2 ;
  RECT 264.640 4.600 264.800 4.700 ;
  LAYER ME1 ;
  RECT 264.640 4.600 264.800 4.700 ;
  LAYER VI1 ;
  RECT 264.670 4.600 264.770 4.700 ;
  LAYER VI2 ;
  RECT 264.670 4.600 264.770 4.700 ;
  LAYER VI3 ;
  RECT 264.670 4.600 264.770 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[114]
PIN DI[113]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 261.140 4.600 261.300 4.700 ;
  LAYER ME2 ;
  RECT 261.140 4.600 261.300 4.700 ;
  LAYER ME1 ;
  RECT 261.140 4.600 261.300 4.700 ;
  LAYER VI1 ;
  RECT 261.170 4.600 261.270 4.700 ;
  LAYER VI2 ;
  RECT 261.170 4.600 261.270 4.700 ;
  LAYER VI3 ;
  RECT 261.170 4.600 261.270 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[113]
PIN DO[113]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 262.540 4.600 262.700 4.700 ;
  LAYER ME2 ;
  RECT 262.540 4.600 262.700 4.700 ;
  LAYER ME1 ;
  RECT 262.540 4.600 262.700 4.700 ;
  LAYER VI1 ;
  RECT 262.570 4.600 262.670 4.700 ;
  LAYER VI2 ;
  RECT 262.570 4.600 262.670 4.700 ;
  LAYER VI3 ;
  RECT 262.570 4.600 262.670 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[113]
PIN DI[112]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 259.040 4.600 259.200 4.700 ;
  LAYER ME2 ;
  RECT 259.040 4.600 259.200 4.700 ;
  LAYER ME1 ;
  RECT 259.040 4.600 259.200 4.700 ;
  LAYER VI1 ;
  RECT 259.070 4.600 259.170 4.700 ;
  LAYER VI2 ;
  RECT 259.070 4.600 259.170 4.700 ;
  LAYER VI3 ;
  RECT 259.070 4.600 259.170 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[112]
PIN DO[112]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 260.440 4.600 260.600 4.700 ;
  LAYER ME2 ;
  RECT 260.440 4.600 260.600 4.700 ;
  LAYER ME1 ;
  RECT 260.440 4.600 260.600 4.700 ;
  LAYER VI1 ;
  RECT 260.470 4.600 260.570 4.700 ;
  LAYER VI2 ;
  RECT 260.470 4.600 260.570 4.700 ;
  LAYER VI3 ;
  RECT 260.470 4.600 260.570 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[112]
PIN DI[111]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 256.940 4.600 257.100 4.700 ;
  LAYER ME2 ;
  RECT 256.940 4.600 257.100 4.700 ;
  LAYER ME1 ;
  RECT 256.940 4.600 257.100 4.700 ;
  LAYER VI1 ;
  RECT 256.970 4.600 257.070 4.700 ;
  LAYER VI2 ;
  RECT 256.970 4.600 257.070 4.700 ;
  LAYER VI3 ;
  RECT 256.970 4.600 257.070 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[111]
PIN DO[111]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 258.340 4.600 258.500 4.700 ;
  LAYER ME2 ;
  RECT 258.340 4.600 258.500 4.700 ;
  LAYER ME1 ;
  RECT 258.340 4.600 258.500 4.700 ;
  LAYER VI1 ;
  RECT 258.370 4.600 258.470 4.700 ;
  LAYER VI2 ;
  RECT 258.370 4.600 258.470 4.700 ;
  LAYER VI3 ;
  RECT 258.370 4.600 258.470 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[111]
PIN DI[110]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 254.840 4.600 255.000 4.700 ;
  LAYER ME2 ;
  RECT 254.840 4.600 255.000 4.700 ;
  LAYER ME1 ;
  RECT 254.840 4.600 255.000 4.700 ;
  LAYER VI1 ;
  RECT 254.870 4.600 254.970 4.700 ;
  LAYER VI2 ;
  RECT 254.870 4.600 254.970 4.700 ;
  LAYER VI3 ;
  RECT 254.870 4.600 254.970 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[110]
PIN DO[110]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 256.240 4.600 256.400 4.700 ;
  LAYER ME2 ;
  RECT 256.240 4.600 256.400 4.700 ;
  LAYER ME1 ;
  RECT 256.240 4.600 256.400 4.700 ;
  LAYER VI1 ;
  RECT 256.270 4.600 256.370 4.700 ;
  LAYER VI2 ;
  RECT 256.270 4.600 256.370 4.700 ;
  LAYER VI3 ;
  RECT 256.270 4.600 256.370 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[110]
PIN DI[109]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 252.740 4.600 252.900 4.700 ;
  LAYER ME2 ;
  RECT 252.740 4.600 252.900 4.700 ;
  LAYER ME1 ;
  RECT 252.740 4.600 252.900 4.700 ;
  LAYER VI1 ;
  RECT 252.770 4.600 252.870 4.700 ;
  LAYER VI2 ;
  RECT 252.770 4.600 252.870 4.700 ;
  LAYER VI3 ;
  RECT 252.770 4.600 252.870 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[109]
PIN DO[109]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 254.140 4.600 254.300 4.700 ;
  LAYER ME2 ;
  RECT 254.140 4.600 254.300 4.700 ;
  LAYER ME1 ;
  RECT 254.140 4.600 254.300 4.700 ;
  LAYER VI1 ;
  RECT 254.170 4.600 254.270 4.700 ;
  LAYER VI2 ;
  RECT 254.170 4.600 254.270 4.700 ;
  LAYER VI3 ;
  RECT 254.170 4.600 254.270 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[109]
PIN DI[108]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 250.640 4.600 250.800 4.700 ;
  LAYER ME2 ;
  RECT 250.640 4.600 250.800 4.700 ;
  LAYER ME1 ;
  RECT 250.640 4.600 250.800 4.700 ;
  LAYER VI1 ;
  RECT 250.670 4.600 250.770 4.700 ;
  LAYER VI2 ;
  RECT 250.670 4.600 250.770 4.700 ;
  LAYER VI3 ;
  RECT 250.670 4.600 250.770 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[108]
PIN DO[108]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 252.040 4.600 252.200 4.700 ;
  LAYER ME2 ;
  RECT 252.040 4.600 252.200 4.700 ;
  LAYER ME1 ;
  RECT 252.040 4.600 252.200 4.700 ;
  LAYER VI1 ;
  RECT 252.070 4.600 252.170 4.700 ;
  LAYER VI2 ;
  RECT 252.070 4.600 252.170 4.700 ;
  LAYER VI3 ;
  RECT 252.070 4.600 252.170 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[108]
PIN DI[107]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 248.540 4.600 248.700 4.700 ;
  LAYER ME2 ;
  RECT 248.540 4.600 248.700 4.700 ;
  LAYER ME1 ;
  RECT 248.540 4.600 248.700 4.700 ;
  LAYER VI1 ;
  RECT 248.570 4.600 248.670 4.700 ;
  LAYER VI2 ;
  RECT 248.570 4.600 248.670 4.700 ;
  LAYER VI3 ;
  RECT 248.570 4.600 248.670 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[107]
PIN DO[107]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 249.940 4.600 250.100 4.700 ;
  LAYER ME2 ;
  RECT 249.940 4.600 250.100 4.700 ;
  LAYER ME1 ;
  RECT 249.940 4.600 250.100 4.700 ;
  LAYER VI1 ;
  RECT 249.970 4.600 250.070 4.700 ;
  LAYER VI2 ;
  RECT 249.970 4.600 250.070 4.700 ;
  LAYER VI3 ;
  RECT 249.970 4.600 250.070 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[107]
PIN DI[106]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 246.440 4.600 246.600 4.700 ;
  LAYER ME2 ;
  RECT 246.440 4.600 246.600 4.700 ;
  LAYER ME1 ;
  RECT 246.440 4.600 246.600 4.700 ;
  LAYER VI1 ;
  RECT 246.470 4.600 246.570 4.700 ;
  LAYER VI2 ;
  RECT 246.470 4.600 246.570 4.700 ;
  LAYER VI3 ;
  RECT 246.470 4.600 246.570 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[106]
PIN DO[106]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 247.840 4.600 248.000 4.700 ;
  LAYER ME2 ;
  RECT 247.840 4.600 248.000 4.700 ;
  LAYER ME1 ;
  RECT 247.840 4.600 248.000 4.700 ;
  LAYER VI1 ;
  RECT 247.870 4.600 247.970 4.700 ;
  LAYER VI2 ;
  RECT 247.870 4.600 247.970 4.700 ;
  LAYER VI3 ;
  RECT 247.870 4.600 247.970 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[106]
PIN DI[105]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 244.340 4.600 244.500 4.700 ;
  LAYER ME2 ;
  RECT 244.340 4.600 244.500 4.700 ;
  LAYER ME1 ;
  RECT 244.340 4.600 244.500 4.700 ;
  LAYER VI1 ;
  RECT 244.370 4.600 244.470 4.700 ;
  LAYER VI2 ;
  RECT 244.370 4.600 244.470 4.700 ;
  LAYER VI3 ;
  RECT 244.370 4.600 244.470 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[105]
PIN DO[105]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 245.740 4.600 245.900 4.700 ;
  LAYER ME2 ;
  RECT 245.740 4.600 245.900 4.700 ;
  LAYER ME1 ;
  RECT 245.740 4.600 245.900 4.700 ;
  LAYER VI1 ;
  RECT 245.770 4.600 245.870 4.700 ;
  LAYER VI2 ;
  RECT 245.770 4.600 245.870 4.700 ;
  LAYER VI3 ;
  RECT 245.770 4.600 245.870 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[105]
PIN DI[104]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 242.240 4.600 242.400 4.700 ;
  LAYER ME2 ;
  RECT 242.240 4.600 242.400 4.700 ;
  LAYER ME1 ;
  RECT 242.240 4.600 242.400 4.700 ;
  LAYER VI1 ;
  RECT 242.270 4.600 242.370 4.700 ;
  LAYER VI2 ;
  RECT 242.270 4.600 242.370 4.700 ;
  LAYER VI3 ;
  RECT 242.270 4.600 242.370 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[104]
PIN DO[104]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 243.640 4.600 243.800 4.700 ;
  LAYER ME2 ;
  RECT 243.640 4.600 243.800 4.700 ;
  LAYER ME1 ;
  RECT 243.640 4.600 243.800 4.700 ;
  LAYER VI1 ;
  RECT 243.670 4.600 243.770 4.700 ;
  LAYER VI2 ;
  RECT 243.670 4.600 243.770 4.700 ;
  LAYER VI3 ;
  RECT 243.670 4.600 243.770 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[104]
PIN DI[103]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 240.140 4.600 240.300 4.700 ;
  LAYER ME2 ;
  RECT 240.140 4.600 240.300 4.700 ;
  LAYER ME1 ;
  RECT 240.140 4.600 240.300 4.700 ;
  LAYER VI1 ;
  RECT 240.170 4.600 240.270 4.700 ;
  LAYER VI2 ;
  RECT 240.170 4.600 240.270 4.700 ;
  LAYER VI3 ;
  RECT 240.170 4.600 240.270 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[103]
PIN DO[103]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 241.540 4.600 241.700 4.700 ;
  LAYER ME2 ;
  RECT 241.540 4.600 241.700 4.700 ;
  LAYER ME1 ;
  RECT 241.540 4.600 241.700 4.700 ;
  LAYER VI1 ;
  RECT 241.570 4.600 241.670 4.700 ;
  LAYER VI2 ;
  RECT 241.570 4.600 241.670 4.700 ;
  LAYER VI3 ;
  RECT 241.570 4.600 241.670 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[103]
PIN DI[102]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 238.040 4.600 238.200 4.700 ;
  LAYER ME2 ;
  RECT 238.040 4.600 238.200 4.700 ;
  LAYER ME1 ;
  RECT 238.040 4.600 238.200 4.700 ;
  LAYER VI1 ;
  RECT 238.070 4.600 238.170 4.700 ;
  LAYER VI2 ;
  RECT 238.070 4.600 238.170 4.700 ;
  LAYER VI3 ;
  RECT 238.070 4.600 238.170 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[102]
PIN DO[102]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 239.440 4.600 239.600 4.700 ;
  LAYER ME2 ;
  RECT 239.440 4.600 239.600 4.700 ;
  LAYER ME1 ;
  RECT 239.440 4.600 239.600 4.700 ;
  LAYER VI1 ;
  RECT 239.470 4.600 239.570 4.700 ;
  LAYER VI2 ;
  RECT 239.470 4.600 239.570 4.700 ;
  LAYER VI3 ;
  RECT 239.470 4.600 239.570 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[102]
PIN DI[101]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 235.940 4.600 236.100 4.700 ;
  LAYER ME2 ;
  RECT 235.940 4.600 236.100 4.700 ;
  LAYER ME1 ;
  RECT 235.940 4.600 236.100 4.700 ;
  LAYER VI1 ;
  RECT 235.970 4.600 236.070 4.700 ;
  LAYER VI2 ;
  RECT 235.970 4.600 236.070 4.700 ;
  LAYER VI3 ;
  RECT 235.970 4.600 236.070 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[101]
PIN DO[101]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 237.340 4.600 237.500 4.700 ;
  LAYER ME2 ;
  RECT 237.340 4.600 237.500 4.700 ;
  LAYER ME1 ;
  RECT 237.340 4.600 237.500 4.700 ;
  LAYER VI1 ;
  RECT 237.370 4.600 237.470 4.700 ;
  LAYER VI2 ;
  RECT 237.370 4.600 237.470 4.700 ;
  LAYER VI3 ;
  RECT 237.370 4.600 237.470 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[101]
PIN DI[100]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 233.840 4.600 234.000 4.700 ;
  LAYER ME2 ;
  RECT 233.840 4.600 234.000 4.700 ;
  LAYER ME1 ;
  RECT 233.840 4.600 234.000 4.700 ;
  LAYER VI1 ;
  RECT 233.870 4.600 233.970 4.700 ;
  LAYER VI2 ;
  RECT 233.870 4.600 233.970 4.700 ;
  LAYER VI3 ;
  RECT 233.870 4.600 233.970 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[100]
PIN DO[100]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 235.240 4.600 235.400 4.700 ;
  LAYER ME2 ;
  RECT 235.240 4.600 235.400 4.700 ;
  LAYER ME1 ;
  RECT 235.240 4.600 235.400 4.700 ;
  LAYER VI1 ;
  RECT 235.270 4.600 235.370 4.700 ;
  LAYER VI2 ;
  RECT 235.270 4.600 235.370 4.700 ;
  LAYER VI3 ;
  RECT 235.270 4.600 235.370 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[100]
PIN DI[99]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 231.740 4.600 231.900 4.700 ;
  LAYER ME2 ;
  RECT 231.740 4.600 231.900 4.700 ;
  LAYER ME1 ;
  RECT 231.740 4.600 231.900 4.700 ;
  LAYER VI1 ;
  RECT 231.770 4.600 231.870 4.700 ;
  LAYER VI2 ;
  RECT 231.770 4.600 231.870 4.700 ;
  LAYER VI3 ;
  RECT 231.770 4.600 231.870 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[99]
PIN DO[99]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 233.140 4.600 233.300 4.700 ;
  LAYER ME2 ;
  RECT 233.140 4.600 233.300 4.700 ;
  LAYER ME1 ;
  RECT 233.140 4.600 233.300 4.700 ;
  LAYER VI1 ;
  RECT 233.170 4.600 233.270 4.700 ;
  LAYER VI2 ;
  RECT 233.170 4.600 233.270 4.700 ;
  LAYER VI3 ;
  RECT 233.170 4.600 233.270 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[99]
PIN DI[98]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 229.640 4.600 229.800 4.700 ;
  LAYER ME2 ;
  RECT 229.640 4.600 229.800 4.700 ;
  LAYER ME1 ;
  RECT 229.640 4.600 229.800 4.700 ;
  LAYER VI1 ;
  RECT 229.670 4.600 229.770 4.700 ;
  LAYER VI2 ;
  RECT 229.670 4.600 229.770 4.700 ;
  LAYER VI3 ;
  RECT 229.670 4.600 229.770 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[98]
PIN DO[98]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 231.040 4.600 231.200 4.700 ;
  LAYER ME2 ;
  RECT 231.040 4.600 231.200 4.700 ;
  LAYER ME1 ;
  RECT 231.040 4.600 231.200 4.700 ;
  LAYER VI1 ;
  RECT 231.070 4.600 231.170 4.700 ;
  LAYER VI2 ;
  RECT 231.070 4.600 231.170 4.700 ;
  LAYER VI3 ;
  RECT 231.070 4.600 231.170 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[98]
PIN DI[97]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 227.540 4.600 227.700 4.700 ;
  LAYER ME2 ;
  RECT 227.540 4.600 227.700 4.700 ;
  LAYER ME1 ;
  RECT 227.540 4.600 227.700 4.700 ;
  LAYER VI1 ;
  RECT 227.570 4.600 227.670 4.700 ;
  LAYER VI2 ;
  RECT 227.570 4.600 227.670 4.700 ;
  LAYER VI3 ;
  RECT 227.570 4.600 227.670 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[97]
PIN DO[97]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 228.940 4.600 229.100 4.700 ;
  LAYER ME2 ;
  RECT 228.940 4.600 229.100 4.700 ;
  LAYER ME1 ;
  RECT 228.940 4.600 229.100 4.700 ;
  LAYER VI1 ;
  RECT 228.970 4.600 229.070 4.700 ;
  LAYER VI2 ;
  RECT 228.970 4.600 229.070 4.700 ;
  LAYER VI3 ;
  RECT 228.970 4.600 229.070 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[97]
PIN DI[96]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 225.440 4.600 225.600 4.700 ;
  LAYER ME2 ;
  RECT 225.440 4.600 225.600 4.700 ;
  LAYER ME1 ;
  RECT 225.440 4.600 225.600 4.700 ;
  LAYER VI1 ;
  RECT 225.470 4.600 225.570 4.700 ;
  LAYER VI2 ;
  RECT 225.470 4.600 225.570 4.700 ;
  LAYER VI3 ;
  RECT 225.470 4.600 225.570 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.088 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.464 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       25.188 LAYER ME2 ;
 ANTENNAMAXAREACAR                       27.726 LAYER ME3 ;
END DI[96]
PIN DO[96]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 226.840 4.600 227.000 4.700 ;
  LAYER ME2 ;
  RECT 226.840 4.600 227.000 4.700 ;
  LAYER ME1 ;
  RECT 226.840 4.600 227.000 4.700 ;
  LAYER VI1 ;
  RECT 226.870 4.600 226.970 4.700 ;
  LAYER VI2 ;
  RECT 226.870 4.600 226.970 4.700 ;
  LAYER VI3 ;
  RECT 226.870 4.600 226.970 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[96]
PIN WEB[3]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 225.710 4.600 225.870 4.700 ;
  LAYER ME2 ;
  RECT 225.710 4.600 225.870 4.700 ;
  LAYER ME1 ;
  RECT 225.710 4.600 225.870 4.700 ;
  LAYER VI1 ;
  RECT 225.740 4.600 225.840 4.700 ;
  LAYER VI2 ;
  RECT 225.740 4.600 225.840 4.700 ;
  LAYER VI3 ;
  RECT 225.740 4.600 225.840 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.093 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.124 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.588 LAYER ME2 ;
 ANTENNAGATEAREA                          0.588 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                        0.618 LAYER ME2 ;
 ANTENNAMAXAREACAR                        0.708 LAYER ME3 ;
END WEB[3]
PIN DI[95]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 223.340 4.600 223.500 4.700 ;
  LAYER ME2 ;
  RECT 223.340 4.600 223.500 4.700 ;
  LAYER ME1 ;
  RECT 223.340 4.600 223.500 4.700 ;
  LAYER VI1 ;
  RECT 223.370 4.600 223.470 4.700 ;
  LAYER VI2 ;
  RECT 223.370 4.600 223.470 4.700 ;
  LAYER VI3 ;
  RECT 223.370 4.600 223.470 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[95]
PIN DO[95]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 224.740 4.600 224.900 4.700 ;
  LAYER ME2 ;
  RECT 224.740 4.600 224.900 4.700 ;
  LAYER ME1 ;
  RECT 224.740 4.600 224.900 4.700 ;
  LAYER VI1 ;
  RECT 224.770 4.600 224.870 4.700 ;
  LAYER VI2 ;
  RECT 224.770 4.600 224.870 4.700 ;
  LAYER VI3 ;
  RECT 224.770 4.600 224.870 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[95]
PIN DI[94]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 221.240 4.600 221.400 4.700 ;
  LAYER ME2 ;
  RECT 221.240 4.600 221.400 4.700 ;
  LAYER ME1 ;
  RECT 221.240 4.600 221.400 4.700 ;
  LAYER VI1 ;
  RECT 221.270 4.600 221.370 4.700 ;
  LAYER VI2 ;
  RECT 221.270 4.600 221.370 4.700 ;
  LAYER VI3 ;
  RECT 221.270 4.600 221.370 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[94]
PIN DO[94]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 222.640 4.600 222.800 4.700 ;
  LAYER ME2 ;
  RECT 222.640 4.600 222.800 4.700 ;
  LAYER ME1 ;
  RECT 222.640 4.600 222.800 4.700 ;
  LAYER VI1 ;
  RECT 222.670 4.600 222.770 4.700 ;
  LAYER VI2 ;
  RECT 222.670 4.600 222.770 4.700 ;
  LAYER VI3 ;
  RECT 222.670 4.600 222.770 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[94]
PIN DI[93]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 219.140 4.600 219.300 4.700 ;
  LAYER ME2 ;
  RECT 219.140 4.600 219.300 4.700 ;
  LAYER ME1 ;
  RECT 219.140 4.600 219.300 4.700 ;
  LAYER VI1 ;
  RECT 219.170 4.600 219.270 4.700 ;
  LAYER VI2 ;
  RECT 219.170 4.600 219.270 4.700 ;
  LAYER VI3 ;
  RECT 219.170 4.600 219.270 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[93]
PIN DO[93]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 220.540 4.600 220.700 4.700 ;
  LAYER ME2 ;
  RECT 220.540 4.600 220.700 4.700 ;
  LAYER ME1 ;
  RECT 220.540 4.600 220.700 4.700 ;
  LAYER VI1 ;
  RECT 220.570 4.600 220.670 4.700 ;
  LAYER VI2 ;
  RECT 220.570 4.600 220.670 4.700 ;
  LAYER VI3 ;
  RECT 220.570 4.600 220.670 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[93]
PIN DI[92]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 217.040 4.600 217.200 4.700 ;
  LAYER ME2 ;
  RECT 217.040 4.600 217.200 4.700 ;
  LAYER ME1 ;
  RECT 217.040 4.600 217.200 4.700 ;
  LAYER VI1 ;
  RECT 217.070 4.600 217.170 4.700 ;
  LAYER VI2 ;
  RECT 217.070 4.600 217.170 4.700 ;
  LAYER VI3 ;
  RECT 217.070 4.600 217.170 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[92]
PIN DO[92]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 218.440 4.600 218.600 4.700 ;
  LAYER ME2 ;
  RECT 218.440 4.600 218.600 4.700 ;
  LAYER ME1 ;
  RECT 218.440 4.600 218.600 4.700 ;
  LAYER VI1 ;
  RECT 218.470 4.600 218.570 4.700 ;
  LAYER VI2 ;
  RECT 218.470 4.600 218.570 4.700 ;
  LAYER VI3 ;
  RECT 218.470 4.600 218.570 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[92]
PIN DI[91]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 214.940 4.600 215.100 4.700 ;
  LAYER ME2 ;
  RECT 214.940 4.600 215.100 4.700 ;
  LAYER ME1 ;
  RECT 214.940 4.600 215.100 4.700 ;
  LAYER VI1 ;
  RECT 214.970 4.600 215.070 4.700 ;
  LAYER VI2 ;
  RECT 214.970 4.600 215.070 4.700 ;
  LAYER VI3 ;
  RECT 214.970 4.600 215.070 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[91]
PIN DO[91]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 216.340 4.600 216.500 4.700 ;
  LAYER ME2 ;
  RECT 216.340 4.600 216.500 4.700 ;
  LAYER ME1 ;
  RECT 216.340 4.600 216.500 4.700 ;
  LAYER VI1 ;
  RECT 216.370 4.600 216.470 4.700 ;
  LAYER VI2 ;
  RECT 216.370 4.600 216.470 4.700 ;
  LAYER VI3 ;
  RECT 216.370 4.600 216.470 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[91]
PIN DI[90]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 212.840 4.600 213.000 4.700 ;
  LAYER ME2 ;
  RECT 212.840 4.600 213.000 4.700 ;
  LAYER ME1 ;
  RECT 212.840 4.600 213.000 4.700 ;
  LAYER VI1 ;
  RECT 212.870 4.600 212.970 4.700 ;
  LAYER VI2 ;
  RECT 212.870 4.600 212.970 4.700 ;
  LAYER VI3 ;
  RECT 212.870 4.600 212.970 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[90]
PIN DO[90]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 214.240 4.600 214.400 4.700 ;
  LAYER ME2 ;
  RECT 214.240 4.600 214.400 4.700 ;
  LAYER ME1 ;
  RECT 214.240 4.600 214.400 4.700 ;
  LAYER VI1 ;
  RECT 214.270 4.600 214.370 4.700 ;
  LAYER VI2 ;
  RECT 214.270 4.600 214.370 4.700 ;
  LAYER VI3 ;
  RECT 214.270 4.600 214.370 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[90]
PIN DI[89]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 210.740 4.600 210.900 4.700 ;
  LAYER ME2 ;
  RECT 210.740 4.600 210.900 4.700 ;
  LAYER ME1 ;
  RECT 210.740 4.600 210.900 4.700 ;
  LAYER VI1 ;
  RECT 210.770 4.600 210.870 4.700 ;
  LAYER VI2 ;
  RECT 210.770 4.600 210.870 4.700 ;
  LAYER VI3 ;
  RECT 210.770 4.600 210.870 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[89]
PIN DO[89]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 212.140 4.600 212.300 4.700 ;
  LAYER ME2 ;
  RECT 212.140 4.600 212.300 4.700 ;
  LAYER ME1 ;
  RECT 212.140 4.600 212.300 4.700 ;
  LAYER VI1 ;
  RECT 212.170 4.600 212.270 4.700 ;
  LAYER VI2 ;
  RECT 212.170 4.600 212.270 4.700 ;
  LAYER VI3 ;
  RECT 212.170 4.600 212.270 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[89]
PIN DI[88]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 208.640 4.600 208.800 4.700 ;
  LAYER ME2 ;
  RECT 208.640 4.600 208.800 4.700 ;
  LAYER ME1 ;
  RECT 208.640 4.600 208.800 4.700 ;
  LAYER VI1 ;
  RECT 208.670 4.600 208.770 4.700 ;
  LAYER VI2 ;
  RECT 208.670 4.600 208.770 4.700 ;
  LAYER VI3 ;
  RECT 208.670 4.600 208.770 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[88]
PIN DO[88]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 210.040 4.600 210.200 4.700 ;
  LAYER ME2 ;
  RECT 210.040 4.600 210.200 4.700 ;
  LAYER ME1 ;
  RECT 210.040 4.600 210.200 4.700 ;
  LAYER VI1 ;
  RECT 210.070 4.600 210.170 4.700 ;
  LAYER VI2 ;
  RECT 210.070 4.600 210.170 4.700 ;
  LAYER VI3 ;
  RECT 210.070 4.600 210.170 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[88]
PIN DI[87]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 206.540 4.600 206.700 4.700 ;
  LAYER ME2 ;
  RECT 206.540 4.600 206.700 4.700 ;
  LAYER ME1 ;
  RECT 206.540 4.600 206.700 4.700 ;
  LAYER VI1 ;
  RECT 206.570 4.600 206.670 4.700 ;
  LAYER VI2 ;
  RECT 206.570 4.600 206.670 4.700 ;
  LAYER VI3 ;
  RECT 206.570 4.600 206.670 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[87]
PIN DO[87]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 207.940 4.600 208.100 4.700 ;
  LAYER ME2 ;
  RECT 207.940 4.600 208.100 4.700 ;
  LAYER ME1 ;
  RECT 207.940 4.600 208.100 4.700 ;
  LAYER VI1 ;
  RECT 207.970 4.600 208.070 4.700 ;
  LAYER VI2 ;
  RECT 207.970 4.600 208.070 4.700 ;
  LAYER VI3 ;
  RECT 207.970 4.600 208.070 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[87]
PIN DI[86]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 204.440 4.600 204.600 4.700 ;
  LAYER ME2 ;
  RECT 204.440 4.600 204.600 4.700 ;
  LAYER ME1 ;
  RECT 204.440 4.600 204.600 4.700 ;
  LAYER VI1 ;
  RECT 204.470 4.600 204.570 4.700 ;
  LAYER VI2 ;
  RECT 204.470 4.600 204.570 4.700 ;
  LAYER VI3 ;
  RECT 204.470 4.600 204.570 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[86]
PIN DO[86]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 205.840 4.600 206.000 4.700 ;
  LAYER ME2 ;
  RECT 205.840 4.600 206.000 4.700 ;
  LAYER ME1 ;
  RECT 205.840 4.600 206.000 4.700 ;
  LAYER VI1 ;
  RECT 205.870 4.600 205.970 4.700 ;
  LAYER VI2 ;
  RECT 205.870 4.600 205.970 4.700 ;
  LAYER VI3 ;
  RECT 205.870 4.600 205.970 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[86]
PIN DI[85]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 202.340 4.600 202.500 4.700 ;
  LAYER ME2 ;
  RECT 202.340 4.600 202.500 4.700 ;
  LAYER ME1 ;
  RECT 202.340 4.600 202.500 4.700 ;
  LAYER VI1 ;
  RECT 202.370 4.600 202.470 4.700 ;
  LAYER VI2 ;
  RECT 202.370 4.600 202.470 4.700 ;
  LAYER VI3 ;
  RECT 202.370 4.600 202.470 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[85]
PIN DO[85]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 203.740 4.600 203.900 4.700 ;
  LAYER ME2 ;
  RECT 203.740 4.600 203.900 4.700 ;
  LAYER ME1 ;
  RECT 203.740 4.600 203.900 4.700 ;
  LAYER VI1 ;
  RECT 203.770 4.600 203.870 4.700 ;
  LAYER VI2 ;
  RECT 203.770 4.600 203.870 4.700 ;
  LAYER VI3 ;
  RECT 203.770 4.600 203.870 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[85]
PIN DI[84]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 200.240 4.600 200.400 4.700 ;
  LAYER ME2 ;
  RECT 200.240 4.600 200.400 4.700 ;
  LAYER ME1 ;
  RECT 200.240 4.600 200.400 4.700 ;
  LAYER VI1 ;
  RECT 200.270 4.600 200.370 4.700 ;
  LAYER VI2 ;
  RECT 200.270 4.600 200.370 4.700 ;
  LAYER VI3 ;
  RECT 200.270 4.600 200.370 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[84]
PIN DO[84]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 201.640 4.600 201.800 4.700 ;
  LAYER ME2 ;
  RECT 201.640 4.600 201.800 4.700 ;
  LAYER ME1 ;
  RECT 201.640 4.600 201.800 4.700 ;
  LAYER VI1 ;
  RECT 201.670 4.600 201.770 4.700 ;
  LAYER VI2 ;
  RECT 201.670 4.600 201.770 4.700 ;
  LAYER VI3 ;
  RECT 201.670 4.600 201.770 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[84]
PIN DI[83]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 198.140 4.600 198.300 4.700 ;
  LAYER ME2 ;
  RECT 198.140 4.600 198.300 4.700 ;
  LAYER ME1 ;
  RECT 198.140 4.600 198.300 4.700 ;
  LAYER VI1 ;
  RECT 198.170 4.600 198.270 4.700 ;
  LAYER VI2 ;
  RECT 198.170 4.600 198.270 4.700 ;
  LAYER VI3 ;
  RECT 198.170 4.600 198.270 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[83]
PIN DO[83]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 199.540 4.600 199.700 4.700 ;
  LAYER ME2 ;
  RECT 199.540 4.600 199.700 4.700 ;
  LAYER ME1 ;
  RECT 199.540 4.600 199.700 4.700 ;
  LAYER VI1 ;
  RECT 199.570 4.600 199.670 4.700 ;
  LAYER VI2 ;
  RECT 199.570 4.600 199.670 4.700 ;
  LAYER VI3 ;
  RECT 199.570 4.600 199.670 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[83]
PIN DI[82]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 196.040 4.600 196.200 4.700 ;
  LAYER ME2 ;
  RECT 196.040 4.600 196.200 4.700 ;
  LAYER ME1 ;
  RECT 196.040 4.600 196.200 4.700 ;
  LAYER VI1 ;
  RECT 196.070 4.600 196.170 4.700 ;
  LAYER VI2 ;
  RECT 196.070 4.600 196.170 4.700 ;
  LAYER VI3 ;
  RECT 196.070 4.600 196.170 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[82]
PIN DO[82]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 197.440 4.600 197.600 4.700 ;
  LAYER ME2 ;
  RECT 197.440 4.600 197.600 4.700 ;
  LAYER ME1 ;
  RECT 197.440 4.600 197.600 4.700 ;
  LAYER VI1 ;
  RECT 197.470 4.600 197.570 4.700 ;
  LAYER VI2 ;
  RECT 197.470 4.600 197.570 4.700 ;
  LAYER VI3 ;
  RECT 197.470 4.600 197.570 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[82]
PIN DI[81]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 193.940 4.600 194.100 4.700 ;
  LAYER ME2 ;
  RECT 193.940 4.600 194.100 4.700 ;
  LAYER ME1 ;
  RECT 193.940 4.600 194.100 4.700 ;
  LAYER VI1 ;
  RECT 193.970 4.600 194.070 4.700 ;
  LAYER VI2 ;
  RECT 193.970 4.600 194.070 4.700 ;
  LAYER VI3 ;
  RECT 193.970 4.600 194.070 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[81]
PIN DO[81]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 195.340 4.600 195.500 4.700 ;
  LAYER ME2 ;
  RECT 195.340 4.600 195.500 4.700 ;
  LAYER ME1 ;
  RECT 195.340 4.600 195.500 4.700 ;
  LAYER VI1 ;
  RECT 195.370 4.600 195.470 4.700 ;
  LAYER VI2 ;
  RECT 195.370 4.600 195.470 4.700 ;
  LAYER VI3 ;
  RECT 195.370 4.600 195.470 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[81]
PIN DI[80]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 191.840 4.600 192.000 4.700 ;
  LAYER ME2 ;
  RECT 191.840 4.600 192.000 4.700 ;
  LAYER ME1 ;
  RECT 191.840 4.600 192.000 4.700 ;
  LAYER VI1 ;
  RECT 191.870 4.600 191.970 4.700 ;
  LAYER VI2 ;
  RECT 191.870 4.600 191.970 4.700 ;
  LAYER VI3 ;
  RECT 191.870 4.600 191.970 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[80]
PIN DO[80]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 193.240 4.600 193.400 4.700 ;
  LAYER ME2 ;
  RECT 193.240 4.600 193.400 4.700 ;
  LAYER ME1 ;
  RECT 193.240 4.600 193.400 4.700 ;
  LAYER VI1 ;
  RECT 193.270 4.600 193.370 4.700 ;
  LAYER VI2 ;
  RECT 193.270 4.600 193.370 4.700 ;
  LAYER VI3 ;
  RECT 193.270 4.600 193.370 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[80]
PIN DI[79]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 189.740 4.600 189.900 4.700 ;
  LAYER ME2 ;
  RECT 189.740 4.600 189.900 4.700 ;
  LAYER ME1 ;
  RECT 189.740 4.600 189.900 4.700 ;
  LAYER VI1 ;
  RECT 189.770 4.600 189.870 4.700 ;
  LAYER VI2 ;
  RECT 189.770 4.600 189.870 4.700 ;
  LAYER VI3 ;
  RECT 189.770 4.600 189.870 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[79]
PIN DO[79]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 191.140 4.600 191.300 4.700 ;
  LAYER ME2 ;
  RECT 191.140 4.600 191.300 4.700 ;
  LAYER ME1 ;
  RECT 191.140 4.600 191.300 4.700 ;
  LAYER VI1 ;
  RECT 191.170 4.600 191.270 4.700 ;
  LAYER VI2 ;
  RECT 191.170 4.600 191.270 4.700 ;
  LAYER VI3 ;
  RECT 191.170 4.600 191.270 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[79]
PIN DI[78]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 187.640 4.600 187.800 4.700 ;
  LAYER ME2 ;
  RECT 187.640 4.600 187.800 4.700 ;
  LAYER ME1 ;
  RECT 187.640 4.600 187.800 4.700 ;
  LAYER VI1 ;
  RECT 187.670 4.600 187.770 4.700 ;
  LAYER VI2 ;
  RECT 187.670 4.600 187.770 4.700 ;
  LAYER VI3 ;
  RECT 187.670 4.600 187.770 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[78]
PIN DO[78]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 189.040 4.600 189.200 4.700 ;
  LAYER ME2 ;
  RECT 189.040 4.600 189.200 4.700 ;
  LAYER ME1 ;
  RECT 189.040 4.600 189.200 4.700 ;
  LAYER VI1 ;
  RECT 189.070 4.600 189.170 4.700 ;
  LAYER VI2 ;
  RECT 189.070 4.600 189.170 4.700 ;
  LAYER VI3 ;
  RECT 189.070 4.600 189.170 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[78]
PIN DI[77]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 185.540 4.600 185.700 4.700 ;
  LAYER ME2 ;
  RECT 185.540 4.600 185.700 4.700 ;
  LAYER ME1 ;
  RECT 185.540 4.600 185.700 4.700 ;
  LAYER VI1 ;
  RECT 185.570 4.600 185.670 4.700 ;
  LAYER VI2 ;
  RECT 185.570 4.600 185.670 4.700 ;
  LAYER VI3 ;
  RECT 185.570 4.600 185.670 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[77]
PIN DO[77]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 186.940 4.600 187.100 4.700 ;
  LAYER ME2 ;
  RECT 186.940 4.600 187.100 4.700 ;
  LAYER ME1 ;
  RECT 186.940 4.600 187.100 4.700 ;
  LAYER VI1 ;
  RECT 186.970 4.600 187.070 4.700 ;
  LAYER VI2 ;
  RECT 186.970 4.600 187.070 4.700 ;
  LAYER VI3 ;
  RECT 186.970 4.600 187.070 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[77]
PIN DI[76]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 183.440 4.600 183.600 4.700 ;
  LAYER ME2 ;
  RECT 183.440 4.600 183.600 4.700 ;
  LAYER ME1 ;
  RECT 183.440 4.600 183.600 4.700 ;
  LAYER VI1 ;
  RECT 183.470 4.600 183.570 4.700 ;
  LAYER VI2 ;
  RECT 183.470 4.600 183.570 4.700 ;
  LAYER VI3 ;
  RECT 183.470 4.600 183.570 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[76]
PIN DO[76]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 184.840 4.600 185.000 4.700 ;
  LAYER ME2 ;
  RECT 184.840 4.600 185.000 4.700 ;
  LAYER ME1 ;
  RECT 184.840 4.600 185.000 4.700 ;
  LAYER VI1 ;
  RECT 184.870 4.600 184.970 4.700 ;
  LAYER VI2 ;
  RECT 184.870 4.600 184.970 4.700 ;
  LAYER VI3 ;
  RECT 184.870 4.600 184.970 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[76]
PIN DI[75]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 181.340 4.600 181.500 4.700 ;
  LAYER ME2 ;
  RECT 181.340 4.600 181.500 4.700 ;
  LAYER ME1 ;
  RECT 181.340 4.600 181.500 4.700 ;
  LAYER VI1 ;
  RECT 181.370 4.600 181.470 4.700 ;
  LAYER VI2 ;
  RECT 181.370 4.600 181.470 4.700 ;
  LAYER VI3 ;
  RECT 181.370 4.600 181.470 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[75]
PIN DO[75]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 182.740 4.600 182.900 4.700 ;
  LAYER ME2 ;
  RECT 182.740 4.600 182.900 4.700 ;
  LAYER ME1 ;
  RECT 182.740 4.600 182.900 4.700 ;
  LAYER VI1 ;
  RECT 182.770 4.600 182.870 4.700 ;
  LAYER VI2 ;
  RECT 182.770 4.600 182.870 4.700 ;
  LAYER VI3 ;
  RECT 182.770 4.600 182.870 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[75]
PIN DI[74]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 179.240 4.600 179.400 4.700 ;
  LAYER ME2 ;
  RECT 179.240 4.600 179.400 4.700 ;
  LAYER ME1 ;
  RECT 179.240 4.600 179.400 4.700 ;
  LAYER VI1 ;
  RECT 179.270 4.600 179.370 4.700 ;
  LAYER VI2 ;
  RECT 179.270 4.600 179.370 4.700 ;
  LAYER VI3 ;
  RECT 179.270 4.600 179.370 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[74]
PIN DO[74]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 180.640 4.600 180.800 4.700 ;
  LAYER ME2 ;
  RECT 180.640 4.600 180.800 4.700 ;
  LAYER ME1 ;
  RECT 180.640 4.600 180.800 4.700 ;
  LAYER VI1 ;
  RECT 180.670 4.600 180.770 4.700 ;
  LAYER VI2 ;
  RECT 180.670 4.600 180.770 4.700 ;
  LAYER VI3 ;
  RECT 180.670 4.600 180.770 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[74]
PIN DI[73]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 177.140 4.600 177.300 4.700 ;
  LAYER ME2 ;
  RECT 177.140 4.600 177.300 4.700 ;
  LAYER ME1 ;
  RECT 177.140 4.600 177.300 4.700 ;
  LAYER VI1 ;
  RECT 177.170 4.600 177.270 4.700 ;
  LAYER VI2 ;
  RECT 177.170 4.600 177.270 4.700 ;
  LAYER VI3 ;
  RECT 177.170 4.600 177.270 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[73]
PIN DO[73]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 178.540 4.600 178.700 4.700 ;
  LAYER ME2 ;
  RECT 178.540 4.600 178.700 4.700 ;
  LAYER ME1 ;
  RECT 178.540 4.600 178.700 4.700 ;
  LAYER VI1 ;
  RECT 178.570 4.600 178.670 4.700 ;
  LAYER VI2 ;
  RECT 178.570 4.600 178.670 4.700 ;
  LAYER VI3 ;
  RECT 178.570 4.600 178.670 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[73]
PIN DI[72]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 175.040 4.600 175.200 4.700 ;
  LAYER ME2 ;
  RECT 175.040 4.600 175.200 4.700 ;
  LAYER ME1 ;
  RECT 175.040 4.600 175.200 4.700 ;
  LAYER VI1 ;
  RECT 175.070 4.600 175.170 4.700 ;
  LAYER VI2 ;
  RECT 175.070 4.600 175.170 4.700 ;
  LAYER VI3 ;
  RECT 175.070 4.600 175.170 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[72]
PIN DO[72]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 176.440 4.600 176.600 4.700 ;
  LAYER ME2 ;
  RECT 176.440 4.600 176.600 4.700 ;
  LAYER ME1 ;
  RECT 176.440 4.600 176.600 4.700 ;
  LAYER VI1 ;
  RECT 176.470 4.600 176.570 4.700 ;
  LAYER VI2 ;
  RECT 176.470 4.600 176.570 4.700 ;
  LAYER VI3 ;
  RECT 176.470 4.600 176.570 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[72]
PIN DI[71]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 172.940 4.600 173.100 4.700 ;
  LAYER ME2 ;
  RECT 172.940 4.600 173.100 4.700 ;
  LAYER ME1 ;
  RECT 172.940 4.600 173.100 4.700 ;
  LAYER VI1 ;
  RECT 172.970 4.600 173.070 4.700 ;
  LAYER VI2 ;
  RECT 172.970 4.600 173.070 4.700 ;
  LAYER VI3 ;
  RECT 172.970 4.600 173.070 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[71]
PIN DO[71]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 174.340 4.600 174.500 4.700 ;
  LAYER ME2 ;
  RECT 174.340 4.600 174.500 4.700 ;
  LAYER ME1 ;
  RECT 174.340 4.600 174.500 4.700 ;
  LAYER VI1 ;
  RECT 174.370 4.600 174.470 4.700 ;
  LAYER VI2 ;
  RECT 174.370 4.600 174.470 4.700 ;
  LAYER VI3 ;
  RECT 174.370 4.600 174.470 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[71]
PIN DI[70]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 170.840 4.600 171.000 4.700 ;
  LAYER ME2 ;
  RECT 170.840 4.600 171.000 4.700 ;
  LAYER ME1 ;
  RECT 170.840 4.600 171.000 4.700 ;
  LAYER VI1 ;
  RECT 170.870 4.600 170.970 4.700 ;
  LAYER VI2 ;
  RECT 170.870 4.600 170.970 4.700 ;
  LAYER VI3 ;
  RECT 170.870 4.600 170.970 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[70]
PIN DO[70]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 172.240 4.600 172.400 4.700 ;
  LAYER ME2 ;
  RECT 172.240 4.600 172.400 4.700 ;
  LAYER ME1 ;
  RECT 172.240 4.600 172.400 4.700 ;
  LAYER VI1 ;
  RECT 172.270 4.600 172.370 4.700 ;
  LAYER VI2 ;
  RECT 172.270 4.600 172.370 4.700 ;
  LAYER VI3 ;
  RECT 172.270 4.600 172.370 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[70]
PIN DI[69]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 168.740 4.600 168.900 4.700 ;
  LAYER ME2 ;
  RECT 168.740 4.600 168.900 4.700 ;
  LAYER ME1 ;
  RECT 168.740 4.600 168.900 4.700 ;
  LAYER VI1 ;
  RECT 168.770 4.600 168.870 4.700 ;
  LAYER VI2 ;
  RECT 168.770 4.600 168.870 4.700 ;
  LAYER VI3 ;
  RECT 168.770 4.600 168.870 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[69]
PIN DO[69]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 170.140 4.600 170.300 4.700 ;
  LAYER ME2 ;
  RECT 170.140 4.600 170.300 4.700 ;
  LAYER ME1 ;
  RECT 170.140 4.600 170.300 4.700 ;
  LAYER VI1 ;
  RECT 170.170 4.600 170.270 4.700 ;
  LAYER VI2 ;
  RECT 170.170 4.600 170.270 4.700 ;
  LAYER VI3 ;
  RECT 170.170 4.600 170.270 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[69]
PIN DI[68]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 166.640 4.600 166.800 4.700 ;
  LAYER ME2 ;
  RECT 166.640 4.600 166.800 4.700 ;
  LAYER ME1 ;
  RECT 166.640 4.600 166.800 4.700 ;
  LAYER VI1 ;
  RECT 166.670 4.600 166.770 4.700 ;
  LAYER VI2 ;
  RECT 166.670 4.600 166.770 4.700 ;
  LAYER VI3 ;
  RECT 166.670 4.600 166.770 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[68]
PIN DO[68]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 168.040 4.600 168.200 4.700 ;
  LAYER ME2 ;
  RECT 168.040 4.600 168.200 4.700 ;
  LAYER ME1 ;
  RECT 168.040 4.600 168.200 4.700 ;
  LAYER VI1 ;
  RECT 168.070 4.600 168.170 4.700 ;
  LAYER VI2 ;
  RECT 168.070 4.600 168.170 4.700 ;
  LAYER VI3 ;
  RECT 168.070 4.600 168.170 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[68]
PIN DI[67]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 164.540 4.600 164.700 4.700 ;
  LAYER ME2 ;
  RECT 164.540 4.600 164.700 4.700 ;
  LAYER ME1 ;
  RECT 164.540 4.600 164.700 4.700 ;
  LAYER VI1 ;
  RECT 164.570 4.600 164.670 4.700 ;
  LAYER VI2 ;
  RECT 164.570 4.600 164.670 4.700 ;
  LAYER VI3 ;
  RECT 164.570 4.600 164.670 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[67]
PIN DO[67]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 165.940 4.600 166.100 4.700 ;
  LAYER ME2 ;
  RECT 165.940 4.600 166.100 4.700 ;
  LAYER ME1 ;
  RECT 165.940 4.600 166.100 4.700 ;
  LAYER VI1 ;
  RECT 165.970 4.600 166.070 4.700 ;
  LAYER VI2 ;
  RECT 165.970 4.600 166.070 4.700 ;
  LAYER VI3 ;
  RECT 165.970 4.600 166.070 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[67]
PIN DI[66]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 162.440 4.600 162.600 4.700 ;
  LAYER ME2 ;
  RECT 162.440 4.600 162.600 4.700 ;
  LAYER ME1 ;
  RECT 162.440 4.600 162.600 4.700 ;
  LAYER VI1 ;
  RECT 162.470 4.600 162.570 4.700 ;
  LAYER VI2 ;
  RECT 162.470 4.600 162.570 4.700 ;
  LAYER VI3 ;
  RECT 162.470 4.600 162.570 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[66]
PIN DO[66]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 163.840 4.600 164.000 4.700 ;
  LAYER ME2 ;
  RECT 163.840 4.600 164.000 4.700 ;
  LAYER ME1 ;
  RECT 163.840 4.600 164.000 4.700 ;
  LAYER VI1 ;
  RECT 163.870 4.600 163.970 4.700 ;
  LAYER VI2 ;
  RECT 163.870 4.600 163.970 4.700 ;
  LAYER VI3 ;
  RECT 163.870 4.600 163.970 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[66]
PIN DI[65]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 160.340 4.600 160.500 4.700 ;
  LAYER ME2 ;
  RECT 160.340 4.600 160.500 4.700 ;
  LAYER ME1 ;
  RECT 160.340 4.600 160.500 4.700 ;
  LAYER VI1 ;
  RECT 160.370 4.600 160.470 4.700 ;
  LAYER VI2 ;
  RECT 160.370 4.600 160.470 4.700 ;
  LAYER VI3 ;
  RECT 160.370 4.600 160.470 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.063 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.302 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.637 LAYER ME2 ;
 ANTENNAMAXAREACAR                       20.175 LAYER ME3 ;
END DI[65]
PIN DO[65]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 161.740 4.600 161.900 4.700 ;
  LAYER ME2 ;
  RECT 161.740 4.600 161.900 4.700 ;
  LAYER ME1 ;
  RECT 161.740 4.600 161.900 4.700 ;
  LAYER VI1 ;
  RECT 161.770 4.600 161.870 4.700 ;
  LAYER VI2 ;
  RECT 161.770 4.600 161.870 4.700 ;
  LAYER VI3 ;
  RECT 161.770 4.600 161.870 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[65]
PIN DI[64]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 158.240 4.600 158.400 4.700 ;
  LAYER ME2 ;
  RECT 158.240 4.600 158.400 4.700 ;
  LAYER ME1 ;
  RECT 158.240 4.600 158.400 4.700 ;
  LAYER VI1 ;
  RECT 158.270 4.600 158.370 4.700 ;
  LAYER VI2 ;
  RECT 158.270 4.600 158.370 4.700 ;
  LAYER VI3 ;
  RECT 158.270 4.600 158.370 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.088 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.464 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.021 LAYER ME2 ;
 ANTENNAGATEAREA                          0.021 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                       25.188 LAYER ME2 ;
 ANTENNAMAXAREACAR                       27.726 LAYER ME3 ;
END DI[64]
PIN DO[64]
  DIRECTION OUTPUT ;
 PORT
  LAYER ME3 ;
  RECT 159.640 4.600 159.800 4.700 ;
  LAYER ME2 ;
  RECT 159.640 4.600 159.800 4.700 ;
  LAYER ME1 ;
  RECT 159.640 4.600 159.800 4.700 ;
  LAYER VI1 ;
  RECT 159.670 4.600 159.770 4.700 ;
  LAYER VI2 ;
  RECT 159.670 4.600 159.770 4.700 ;
  LAYER VI3 ;
  RECT 159.670 4.600 159.770 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.534 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.252 LAYER ME3 ;
 ANTENNADIFFAREA                          0.594 LAYER ME3 ;
END DO[64]
PIN WEB[2]
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 158.510 4.600 158.670 4.700 ;
  LAYER ME2 ;
  RECT 158.510 4.600 158.670 4.700 ;
  LAYER ME1 ;
  RECT 158.510 4.600 158.670 4.700 ;
  LAYER VI1 ;
  RECT 158.540 4.600 158.640 4.700 ;
  LAYER VI2 ;
  RECT 158.540 4.600 158.640 4.700 ;
  LAYER VI3 ;
  RECT 158.540 4.600 158.640 4.700 ;
 END
 ANTENNAPARTIALMETALAREA                  0.093 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  0.124 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.037 LAYER ME3 ;
 ANTENNAGATEAREA                          0.588 LAYER ME2 ;
 ANTENNAGATEAREA                          0.588 LAYER ME3 ;
 ANTENNADIFFAREA                          0.058 LAYER ME1 ;
 ANTENNADIFFAREA                          0.058 LAYER ME2 ;
 ANTENNADIFFAREA                          0.058 LAYER ME3 ;
 ANTENNAMAXAREACAR                        0.618 LAYER ME2 ;
 ANTENNAMAXAREACAR                        0.708 LAYER ME3 ;
END WEB[2]
PIN GND
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE RING ;
 PORT
  LAYER ME3 ;
  RECT 0.000 0.000 298.405 2.000 ;
  RECT 0.000 162.840 298.405 164.840 ;
  LAYER ME2 ;
  RECT 296.405 0.000 298.405 164.840 ;
  RECT 0.000 0.000 2.000 164.840 ;
 END
END GND
PIN VCC
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE RING ;
 PORT
  LAYER ME3 ;
  RECT 2.300 2.300 296.105 4.300 ;
  RECT 2.300 160.540 296.105 162.540 ;
  LAYER ME2 ;
  RECT 294.105 2.300 296.105 162.540 ;
  RECT 2.300 2.300 4.300 162.540 ;
 END
END VCC
OBS
  LAYER VI3 SPACING 0.300 ;
  RECT 4.600 4.600 293.805 160.240 ;
  LAYER VI2 SPACING 0.300 ;
  RECT 4.600 4.600 293.805 160.240 ;
  LAYER VI1 SPACING 0.300 ;
  RECT 4.600 4.600 293.805 160.240 ;
  LAYER ME3 SPACING 0.300 ;
  RECT 4.600 4.600 293.805 160.240 ;
  RECT 159.905 2.300 160.215 4.600 ;
  RECT 162.005 2.300 162.315 4.600 ;
  RECT 164.105 2.300 164.415 4.600 ;
  RECT 166.205 2.300 166.515 4.600 ;
  RECT 168.305 2.300 168.615 4.600 ;
  RECT 170.405 2.300 170.715 4.600 ;
  RECT 172.505 2.300 172.815 4.600 ;
  RECT 174.605 2.300 174.915 4.600 ;
  RECT 176.705 2.300 177.015 4.600 ;
  RECT 178.805 2.300 179.115 4.600 ;
  RECT 180.905 2.300 181.215 4.600 ;
  RECT 183.005 2.300 183.315 4.600 ;
  RECT 185.105 2.300 185.415 4.600 ;
  RECT 187.205 2.300 187.515 4.600 ;
  RECT 189.305 2.300 189.615 4.600 ;
  RECT 191.405 2.300 191.715 4.600 ;
  RECT 193.505 2.300 193.815 4.600 ;
  RECT 195.605 2.300 195.915 4.600 ;
  RECT 197.705 2.300 198.015 4.600 ;
  RECT 199.805 2.300 200.115 4.600 ;
  RECT 201.905 2.300 202.215 4.600 ;
  RECT 204.005 2.300 204.315 4.600 ;
  RECT 206.105 2.300 206.415 4.600 ;
  RECT 208.205 2.300 208.515 4.600 ;
  RECT 210.305 2.300 210.615 4.600 ;
  RECT 212.405 2.300 212.715 4.600 ;
  RECT 214.505 2.300 214.815 4.600 ;
  RECT 216.605 2.300 216.915 4.600 ;
  RECT 218.705 2.300 219.015 4.600 ;
  RECT 220.805 2.300 221.115 4.600 ;
  RECT 222.905 2.300 223.215 4.600 ;
  RECT 225.005 2.300 225.315 4.600 ;
  RECT 227.105 2.300 227.415 4.600 ;
  RECT 229.205 2.300 229.515 4.600 ;
  RECT 231.305 2.300 231.615 4.600 ;
  RECT 233.405 2.300 233.715 4.600 ;
  RECT 235.505 2.300 235.815 4.600 ;
  RECT 237.605 2.300 237.915 4.600 ;
  RECT 239.705 2.300 240.015 4.600 ;
  RECT 241.805 2.300 242.115 4.600 ;
  RECT 243.905 2.300 244.215 4.600 ;
  RECT 246.005 2.300 246.315 4.600 ;
  RECT 248.105 2.300 248.415 4.600 ;
  RECT 250.205 2.300 250.515 4.600 ;
  RECT 252.305 2.300 252.615 4.600 ;
  RECT 254.405 2.300 254.715 4.600 ;
  RECT 256.505 2.300 256.815 4.600 ;
  RECT 258.605 2.300 258.915 4.600 ;
  RECT 260.705 2.300 261.015 4.600 ;
  RECT 262.805 2.300 263.115 4.600 ;
  RECT 264.905 2.300 265.215 4.600 ;
  RECT 267.005 2.300 267.315 4.600 ;
  RECT 269.105 2.300 269.415 4.600 ;
  RECT 271.205 2.300 271.515 4.600 ;
  RECT 273.305 2.300 273.615 4.600 ;
  RECT 275.405 2.300 275.715 4.600 ;
  RECT 277.505 2.300 277.815 4.600 ;
  RECT 279.605 2.300 279.915 4.600 ;
  RECT 281.705 2.300 282.015 4.600 ;
  RECT 283.805 2.300 284.115 4.600 ;
  RECT 285.905 2.300 286.215 4.600 ;
  RECT 288.005 2.300 288.315 4.600 ;
  RECT 290.105 2.300 290.415 4.600 ;
  RECT 292.205 2.300 292.515 4.600 ;
  RECT 292.915 2.300 293.225 4.600 ;
  RECT 153.660 2.300 154.180 4.600 ;
  RECT 151.860 2.300 152.380 4.600 ;
  RECT 154.395 2.300 154.915 4.600 ;
  RECT 148.920 2.300 149.400 4.600 ;
  RECT 147.150 2.300 147.530 4.600 ;
  RECT 146.465 2.300 146.775 4.600 ;
  RECT 144.870 2.300 145.250 4.600 ;
  RECT 144.185 2.300 144.495 4.600 ;
  RECT 142.590 2.300 142.970 4.600 ;
  RECT 141.905 2.300 142.215 4.600 ;
  RECT 5.180 2.300 5.490 4.600 ;
  RECT 7.680 2.300 7.990 4.600 ;
  RECT 9.780 2.300 10.090 4.600 ;
  RECT 11.880 2.300 12.190 4.600 ;
  RECT 13.980 2.300 14.290 4.600 ;
  RECT 16.080 2.300 16.390 4.600 ;
  RECT 18.180 2.300 18.490 4.600 ;
  RECT 20.280 2.300 20.590 4.600 ;
  RECT 22.380 2.300 22.690 4.600 ;
  RECT 24.480 2.300 24.790 4.600 ;
  RECT 26.580 2.300 26.890 4.600 ;
  RECT 28.680 2.300 28.990 4.600 ;
  RECT 30.780 2.300 31.090 4.600 ;
  RECT 32.880 2.300 33.190 4.600 ;
  RECT 34.980 2.300 35.290 4.600 ;
  RECT 37.080 2.300 37.390 4.600 ;
  RECT 39.180 2.300 39.490 4.600 ;
  RECT 41.280 2.300 41.590 4.600 ;
  RECT 43.380 2.300 43.690 4.600 ;
  RECT 45.480 2.300 45.790 4.600 ;
  RECT 47.580 2.300 47.890 4.600 ;
  RECT 49.680 2.300 49.990 4.600 ;
  RECT 51.780 2.300 52.090 4.600 ;
  RECT 53.880 2.300 54.190 4.600 ;
  RECT 55.980 2.300 56.290 4.600 ;
  RECT 58.080 2.300 58.390 4.600 ;
  RECT 60.180 2.300 60.490 4.600 ;
  RECT 62.280 2.300 62.590 4.600 ;
  RECT 64.380 2.300 64.690 4.600 ;
  RECT 66.480 2.300 66.790 4.600 ;
  RECT 68.580 2.300 68.890 4.600 ;
  RECT 70.680 2.300 70.990 4.600 ;
  RECT 72.780 2.300 73.090 4.600 ;
  RECT 74.880 2.300 75.190 4.600 ;
  RECT 76.980 2.300 77.290 4.600 ;
  RECT 79.080 2.300 79.390 4.600 ;
  RECT 81.180 2.300 81.490 4.600 ;
  RECT 83.280 2.300 83.590 4.600 ;
  RECT 85.380 2.300 85.690 4.600 ;
  RECT 87.480 2.300 87.790 4.600 ;
  RECT 89.580 2.300 89.890 4.600 ;
  RECT 91.680 2.300 91.990 4.600 ;
  RECT 93.780 2.300 94.090 4.600 ;
  RECT 95.880 2.300 96.190 4.600 ;
  RECT 97.980 2.300 98.290 4.600 ;
  RECT 100.080 2.300 100.390 4.600 ;
  RECT 102.180 2.300 102.490 4.600 ;
  RECT 104.280 2.300 104.590 4.600 ;
  RECT 106.380 2.300 106.690 4.600 ;
  RECT 108.480 2.300 108.790 4.600 ;
  RECT 110.580 2.300 110.890 4.600 ;
  RECT 112.680 2.300 112.990 4.600 ;
  RECT 114.780 2.300 115.090 4.600 ;
  RECT 116.880 2.300 117.190 4.600 ;
  RECT 118.980 2.300 119.290 4.600 ;
  RECT 121.080 2.300 121.390 4.600 ;
  RECT 123.180 2.300 123.490 4.600 ;
  RECT 125.280 2.300 125.590 4.600 ;
  RECT 127.380 2.300 127.690 4.600 ;
  RECT 129.480 2.300 129.790 4.600 ;
  RECT 131.580 2.300 131.890 4.600 ;
  RECT 133.680 2.300 133.990 4.600 ;
  RECT 135.780 2.300 136.090 4.600 ;
  RECT 137.880 2.300 138.190 4.600 ;
  RECT 139.980 2.300 140.290 4.600 ;
  RECT 292.915 160.240 293.225 162.540 ;
  RECT 157.165 160.240 157.475 162.540 ;
  RECT 156.225 160.240 156.535 162.540 ;
  RECT 155.075 160.240 155.595 162.540 ;
  RECT 154.395 160.240 154.915 162.540 ;
  RECT 153.660 160.240 154.180 162.540 ;
  RECT 151.860 160.240 152.380 162.540 ;
  RECT 150.840 160.240 151.150 162.540 ;
  RECT 148.920 160.240 149.400 162.540 ;
  RECT 147.150 160.240 147.530 162.540 ;
  RECT 144.185 160.240 144.495 162.540 ;
  RECT 142.590 160.240 142.970 162.540 ;
  RECT 141.905 160.240 142.215 162.540 ;
  RECT 146.465 160.240 146.775 162.540 ;
  RECT 144.870 160.240 145.250 162.540 ;
  RECT 5.180 160.240 5.490 162.540 ;
  RECT 140.560 160.240 140.710 162.540 ;
  RECT 0.000 0.000 298.405 2.000 ;
  RECT 0.000 162.840 298.405 164.840 ;
  RECT 2.300 2.300 296.105 4.300 ;
  RECT 2.300 160.540 296.105 162.540 ;
  LAYER ME2 SPACING 0.300 ;
  RECT 4.600 4.600 293.805 160.240 ;
  RECT 159.220 0.000 159.530 4.600 ;
  RECT 158.770 0.000 159.080 4.600 ;
  RECT 160.870 0.000 161.180 4.600 ;
  RECT 161.320 0.000 161.630 4.600 ;
  RECT 162.970 0.000 163.280 4.600 ;
  RECT 163.420 0.000 163.730 4.600 ;
  RECT 165.070 0.000 165.380 4.600 ;
  RECT 165.520 0.000 165.830 4.600 ;
  RECT 167.170 0.000 167.480 4.600 ;
  RECT 167.620 0.000 167.930 4.600 ;
  RECT 169.270 0.000 169.580 4.600 ;
  RECT 169.720 0.000 170.030 4.600 ;
  RECT 171.370 0.000 171.680 4.600 ;
  RECT 171.820 0.000 172.130 4.600 ;
  RECT 173.470 0.000 173.780 4.600 ;
  RECT 173.920 0.000 174.230 4.600 ;
  RECT 175.570 0.000 175.880 4.600 ;
  RECT 176.020 0.000 176.330 4.600 ;
  RECT 177.670 0.000 177.980 4.600 ;
  RECT 178.120 0.000 178.430 4.600 ;
  RECT 179.770 0.000 180.080 4.600 ;
  RECT 180.220 0.000 180.530 4.600 ;
  RECT 181.870 0.000 182.180 4.600 ;
  RECT 182.320 0.000 182.630 4.600 ;
  RECT 183.970 0.000 184.280 4.600 ;
  RECT 184.420 0.000 184.730 4.600 ;
  RECT 186.070 0.000 186.380 4.600 ;
  RECT 186.520 0.000 186.830 4.600 ;
  RECT 188.170 0.000 188.480 4.600 ;
  RECT 188.620 0.000 188.930 4.600 ;
  RECT 190.270 0.000 190.580 4.600 ;
  RECT 190.720 0.000 191.030 4.600 ;
  RECT 192.370 0.000 192.680 4.600 ;
  RECT 192.820 0.000 193.130 4.600 ;
  RECT 194.470 0.000 194.780 4.600 ;
  RECT 194.920 0.000 195.230 4.600 ;
  RECT 196.570 0.000 196.880 4.600 ;
  RECT 197.020 0.000 197.330 4.600 ;
  RECT 198.670 0.000 198.980 4.600 ;
  RECT 199.120 0.000 199.430 4.600 ;
  RECT 200.770 0.000 201.080 4.600 ;
  RECT 201.220 0.000 201.530 4.600 ;
  RECT 202.870 0.000 203.180 4.600 ;
  RECT 203.320 0.000 203.630 4.600 ;
  RECT 204.970 0.000 205.280 4.600 ;
  RECT 205.420 0.000 205.730 4.600 ;
  RECT 207.070 0.000 207.380 4.600 ;
  RECT 207.520 0.000 207.830 4.600 ;
  RECT 209.170 0.000 209.480 4.600 ;
  RECT 209.620 0.000 209.930 4.600 ;
  RECT 211.270 0.000 211.580 4.600 ;
  RECT 211.720 0.000 212.030 4.600 ;
  RECT 213.370 0.000 213.680 4.600 ;
  RECT 213.820 0.000 214.130 4.600 ;
  RECT 215.470 0.000 215.780 4.600 ;
  RECT 215.920 0.000 216.230 4.600 ;
  RECT 217.570 0.000 217.880 4.600 ;
  RECT 218.020 0.000 218.330 4.600 ;
  RECT 219.670 0.000 219.980 4.600 ;
  RECT 220.120 0.000 220.430 4.600 ;
  RECT 221.770 0.000 222.080 4.600 ;
  RECT 222.220 0.000 222.530 4.600 ;
  RECT 223.870 0.000 224.180 4.600 ;
  RECT 224.320 0.000 224.630 4.600 ;
  RECT 226.420 0.000 226.730 4.600 ;
  RECT 225.970 0.000 226.280 4.600 ;
  RECT 228.070 0.000 228.380 4.600 ;
  RECT 228.520 0.000 228.830 4.600 ;
  RECT 230.170 0.000 230.480 4.600 ;
  RECT 230.620 0.000 230.930 4.600 ;
  RECT 232.270 0.000 232.580 4.600 ;
  RECT 232.720 0.000 233.030 4.600 ;
  RECT 234.370 0.000 234.680 4.600 ;
  RECT 234.820 0.000 235.130 4.600 ;
  RECT 236.470 0.000 236.780 4.600 ;
  RECT 236.920 0.000 237.230 4.600 ;
  RECT 238.570 0.000 238.880 4.600 ;
  RECT 239.020 0.000 239.330 4.600 ;
  RECT 240.670 0.000 240.980 4.600 ;
  RECT 241.120 0.000 241.430 4.600 ;
  RECT 242.770 0.000 243.080 4.600 ;
  RECT 243.220 0.000 243.530 4.600 ;
  RECT 244.870 0.000 245.180 4.600 ;
  RECT 245.320 0.000 245.630 4.600 ;
  RECT 246.970 0.000 247.280 4.600 ;
  RECT 247.420 0.000 247.730 4.600 ;
  RECT 249.070 0.000 249.380 4.600 ;
  RECT 249.520 0.000 249.830 4.600 ;
  RECT 251.170 0.000 251.480 4.600 ;
  RECT 251.620 0.000 251.930 4.600 ;
  RECT 253.270 0.000 253.580 4.600 ;
  RECT 253.720 0.000 254.030 4.600 ;
  RECT 255.370 0.000 255.680 4.600 ;
  RECT 255.820 0.000 256.130 4.600 ;
  RECT 257.470 0.000 257.780 4.600 ;
  RECT 257.920 0.000 258.230 4.600 ;
  RECT 259.570 0.000 259.880 4.600 ;
  RECT 260.020 0.000 260.330 4.600 ;
  RECT 261.670 0.000 261.980 4.600 ;
  RECT 262.120 0.000 262.430 4.600 ;
  RECT 263.770 0.000 264.080 4.600 ;
  RECT 264.220 0.000 264.530 4.600 ;
  RECT 265.870 0.000 266.180 4.600 ;
  RECT 266.320 0.000 266.630 4.600 ;
  RECT 267.970 0.000 268.280 4.600 ;
  RECT 268.420 0.000 268.730 4.600 ;
  RECT 270.070 0.000 270.380 4.600 ;
  RECT 270.520 0.000 270.830 4.600 ;
  RECT 272.170 0.000 272.480 4.600 ;
  RECT 272.620 0.000 272.930 4.600 ;
  RECT 274.270 0.000 274.580 4.600 ;
  RECT 274.720 0.000 275.030 4.600 ;
  RECT 276.370 0.000 276.680 4.600 ;
  RECT 276.820 0.000 277.130 4.600 ;
  RECT 278.470 0.000 278.780 4.600 ;
  RECT 278.920 0.000 279.230 4.600 ;
  RECT 280.570 0.000 280.880 4.600 ;
  RECT 281.020 0.000 281.330 4.600 ;
  RECT 282.670 0.000 282.980 4.600 ;
  RECT 283.120 0.000 283.430 4.600 ;
  RECT 284.770 0.000 285.080 4.600 ;
  RECT 285.220 0.000 285.530 4.600 ;
  RECT 286.870 0.000 287.180 4.600 ;
  RECT 287.320 0.000 287.630 4.600 ;
  RECT 288.970 0.000 289.280 4.600 ;
  RECT 289.420 0.000 289.730 4.600 ;
  RECT 291.070 0.000 291.380 4.600 ;
  RECT 291.520 0.000 291.830 4.600 ;
  RECT 292.645 0.000 292.815 4.600 ;
  RECT 293.805 5.695 296.105 6.215 ;
  RECT 293.805 8.470 296.105 8.990 ;
  RECT 293.805 10.885 296.105 11.195 ;
  RECT 293.805 12.515 296.105 12.825 ;
  RECT 293.805 14.365 296.105 14.885 ;
  RECT 293.805 17.030 296.105 17.550 ;
  RECT 293.805 20.180 296.105 20.700 ;
  RECT 293.805 21.080 296.105 21.390 ;
  RECT 293.805 24.110 296.105 24.420 ;
  RECT 293.805 26.840 296.105 27.420 ;
  RECT 157.750 0.000 158.060 4.600 ;
  RECT 152.690 0.000 153.210 4.600 ;
  RECT 148.050 0.000 148.530 4.600 ;
  RECT 146.055 0.000 146.365 4.600 ;
  RECT 145.380 0.000 145.690 4.600 ;
  RECT 143.775 0.000 144.085 4.600 ;
  RECT 143.100 0.000 143.410 4.600 ;
  RECT 141.495 0.000 141.805 4.600 ;
  RECT 140.820 0.000 141.130 4.600 ;
  RECT 5.590 0.000 5.760 4.600 ;
  RECT 2.300 5.695 4.600 6.215 ;
  RECT 2.300 8.470 4.600 8.990 ;
  RECT 2.300 10.885 4.600 11.195 ;
  RECT 2.300 12.515 4.600 12.825 ;
  RECT 2.300 14.365 4.600 14.885 ;
  RECT 2.300 17.030 4.600 17.550 ;
  RECT 2.300 20.180 4.600 20.700 ;
  RECT 2.300 21.080 4.600 21.390 ;
  RECT 2.300 24.110 4.600 24.420 ;
  RECT 2.300 26.840 4.600 27.420 ;
  RECT 6.995 0.000 7.305 4.600 ;
  RECT 6.545 0.000 6.855 4.600 ;
  RECT 8.645 0.000 8.955 4.600 ;
  RECT 9.095 0.000 9.405 4.600 ;
  RECT 10.745 0.000 11.055 4.600 ;
  RECT 11.195 0.000 11.505 4.600 ;
  RECT 12.845 0.000 13.155 4.600 ;
  RECT 13.295 0.000 13.605 4.600 ;
  RECT 14.945 0.000 15.255 4.600 ;
  RECT 15.395 0.000 15.705 4.600 ;
  RECT 17.045 0.000 17.355 4.600 ;
  RECT 17.495 0.000 17.805 4.600 ;
  RECT 19.145 0.000 19.455 4.600 ;
  RECT 19.595 0.000 19.905 4.600 ;
  RECT 21.245 0.000 21.555 4.600 ;
  RECT 21.695 0.000 22.005 4.600 ;
  RECT 23.345 0.000 23.655 4.600 ;
  RECT 23.795 0.000 24.105 4.600 ;
  RECT 25.445 0.000 25.755 4.600 ;
  RECT 25.895 0.000 26.205 4.600 ;
  RECT 27.545 0.000 27.855 4.600 ;
  RECT 27.995 0.000 28.305 4.600 ;
  RECT 29.645 0.000 29.955 4.600 ;
  RECT 30.095 0.000 30.405 4.600 ;
  RECT 31.745 0.000 32.055 4.600 ;
  RECT 32.195 0.000 32.505 4.600 ;
  RECT 33.845 0.000 34.155 4.600 ;
  RECT 34.295 0.000 34.605 4.600 ;
  RECT 35.945 0.000 36.255 4.600 ;
  RECT 36.395 0.000 36.705 4.600 ;
  RECT 38.045 0.000 38.355 4.600 ;
  RECT 38.495 0.000 38.805 4.600 ;
  RECT 40.145 0.000 40.455 4.600 ;
  RECT 40.595 0.000 40.905 4.600 ;
  RECT 42.245 0.000 42.555 4.600 ;
  RECT 42.695 0.000 43.005 4.600 ;
  RECT 44.345 0.000 44.655 4.600 ;
  RECT 44.795 0.000 45.105 4.600 ;
  RECT 46.445 0.000 46.755 4.600 ;
  RECT 46.895 0.000 47.205 4.600 ;
  RECT 48.545 0.000 48.855 4.600 ;
  RECT 48.995 0.000 49.305 4.600 ;
  RECT 50.645 0.000 50.955 4.600 ;
  RECT 51.095 0.000 51.405 4.600 ;
  RECT 52.745 0.000 53.055 4.600 ;
  RECT 53.195 0.000 53.505 4.600 ;
  RECT 54.845 0.000 55.155 4.600 ;
  RECT 55.295 0.000 55.605 4.600 ;
  RECT 56.945 0.000 57.255 4.600 ;
  RECT 57.395 0.000 57.705 4.600 ;
  RECT 59.045 0.000 59.355 4.600 ;
  RECT 59.495 0.000 59.805 4.600 ;
  RECT 61.145 0.000 61.455 4.600 ;
  RECT 61.595 0.000 61.905 4.600 ;
  RECT 63.245 0.000 63.555 4.600 ;
  RECT 63.695 0.000 64.005 4.600 ;
  RECT 65.345 0.000 65.655 4.600 ;
  RECT 65.795 0.000 66.105 4.600 ;
  RECT 67.445 0.000 67.755 4.600 ;
  RECT 67.895 0.000 68.205 4.600 ;
  RECT 69.545 0.000 69.855 4.600 ;
  RECT 69.995 0.000 70.305 4.600 ;
  RECT 71.645 0.000 71.955 4.600 ;
  RECT 72.095 0.000 72.405 4.600 ;
  RECT 74.195 0.000 74.505 4.600 ;
  RECT 73.745 0.000 74.055 4.600 ;
  RECT 75.845 0.000 76.155 4.600 ;
  RECT 76.295 0.000 76.605 4.600 ;
  RECT 77.945 0.000 78.255 4.600 ;
  RECT 78.395 0.000 78.705 4.600 ;
  RECT 80.045 0.000 80.355 4.600 ;
  RECT 80.495 0.000 80.805 4.600 ;
  RECT 82.145 0.000 82.455 4.600 ;
  RECT 82.595 0.000 82.905 4.600 ;
  RECT 84.245 0.000 84.555 4.600 ;
  RECT 84.695 0.000 85.005 4.600 ;
  RECT 86.345 0.000 86.655 4.600 ;
  RECT 86.795 0.000 87.105 4.600 ;
  RECT 88.445 0.000 88.755 4.600 ;
  RECT 88.895 0.000 89.205 4.600 ;
  RECT 90.545 0.000 90.855 4.600 ;
  RECT 90.995 0.000 91.305 4.600 ;
  RECT 92.645 0.000 92.955 4.600 ;
  RECT 93.095 0.000 93.405 4.600 ;
  RECT 94.745 0.000 95.055 4.600 ;
  RECT 95.195 0.000 95.505 4.600 ;
  RECT 96.845 0.000 97.155 4.600 ;
  RECT 97.295 0.000 97.605 4.600 ;
  RECT 98.945 0.000 99.255 4.600 ;
  RECT 99.395 0.000 99.705 4.600 ;
  RECT 101.045 0.000 101.355 4.600 ;
  RECT 101.495 0.000 101.805 4.600 ;
  RECT 103.145 0.000 103.455 4.600 ;
  RECT 103.595 0.000 103.905 4.600 ;
  RECT 105.245 0.000 105.555 4.600 ;
  RECT 105.695 0.000 106.005 4.600 ;
  RECT 107.345 0.000 107.655 4.600 ;
  RECT 107.795 0.000 108.105 4.600 ;
  RECT 109.445 0.000 109.755 4.600 ;
  RECT 109.895 0.000 110.205 4.600 ;
  RECT 111.545 0.000 111.855 4.600 ;
  RECT 111.995 0.000 112.305 4.600 ;
  RECT 113.645 0.000 113.955 4.600 ;
  RECT 114.095 0.000 114.405 4.600 ;
  RECT 115.745 0.000 116.055 4.600 ;
  RECT 116.195 0.000 116.505 4.600 ;
  RECT 117.845 0.000 118.155 4.600 ;
  RECT 118.295 0.000 118.605 4.600 ;
  RECT 119.945 0.000 120.255 4.600 ;
  RECT 120.395 0.000 120.705 4.600 ;
  RECT 122.045 0.000 122.355 4.600 ;
  RECT 122.495 0.000 122.805 4.600 ;
  RECT 124.145 0.000 124.455 4.600 ;
  RECT 124.595 0.000 124.905 4.600 ;
  RECT 126.245 0.000 126.555 4.600 ;
  RECT 126.695 0.000 127.005 4.600 ;
  RECT 128.345 0.000 128.655 4.600 ;
  RECT 128.795 0.000 129.105 4.600 ;
  RECT 130.445 0.000 130.755 4.600 ;
  RECT 130.895 0.000 131.205 4.600 ;
  RECT 132.545 0.000 132.855 4.600 ;
  RECT 132.995 0.000 133.305 4.600 ;
  RECT 134.645 0.000 134.955 4.600 ;
  RECT 135.095 0.000 135.405 4.600 ;
  RECT 136.745 0.000 137.055 4.600 ;
  RECT 137.195 0.000 137.505 4.600 ;
  RECT 138.845 0.000 139.155 4.600 ;
  RECT 139.295 0.000 139.605 4.600 ;
  RECT 157.750 160.240 158.060 164.840 ;
  RECT 293.805 159.375 296.105 159.515 ;
  RECT 292.645 160.240 292.815 164.840 ;
  RECT 293.805 126.855 296.105 126.995 ;
  RECT 293.805 94.055 296.105 94.195 ;
  RECT 293.805 61.255 296.105 61.395 ;
  RECT 156.695 160.240 157.005 164.840 ;
  RECT 155.755 160.240 156.065 164.840 ;
  RECT 152.690 160.240 153.210 164.840 ;
  RECT 151.310 160.240 151.620 164.840 ;
  RECT 150.285 160.240 150.595 164.840 ;
  RECT 149.765 160.240 150.075 164.840 ;
  RECT 148.050 160.240 148.530 164.840 ;
  RECT 143.775 160.240 144.085 164.840 ;
  RECT 143.100 160.240 143.410 164.840 ;
  RECT 141.495 160.240 141.805 164.840 ;
  RECT 140.870 160.240 141.180 164.840 ;
  RECT 146.055 160.240 146.365 164.840 ;
  RECT 145.380 160.240 145.690 164.840 ;
  RECT 2.300 159.375 4.600 159.515 ;
  RECT 5.590 160.240 5.760 164.840 ;
  RECT 2.300 126.855 4.600 126.995 ;
  RECT 2.300 94.055 4.600 94.195 ;
  RECT 2.300 61.255 4.600 61.395 ;
  RECT 296.405 0.000 298.405 164.840 ;
  RECT 0.000 0.000 2.000 164.840 ;
  RECT 294.105 2.300 296.105 162.540 ;
  RECT 2.300 2.300 4.300 162.540 ;
  LAYER ME1 SPACING 0.300 ;
  RECT 4.600 4.600 293.805 160.240 ;
  RECT 293.805 15.700 298.405 16.010 ;
  RECT 293.805 7.030 298.405 7.340 ;
  RECT 293.805 9.625 298.405 9.935 ;
  RECT 293.805 11.415 298.405 11.725 ;
  RECT 293.805 13.465 298.405 13.775 ;
  RECT 293.805 17.845 298.405 18.345 ;
  RECT 293.805 22.535 298.405 22.845 ;
  RECT 293.805 21.590 298.405 21.900 ;
  RECT 293.805 23.700 298.405 24.010 ;
  RECT 293.805 25.860 298.405 26.230 ;
  RECT 0.000 7.030 4.600 7.340 ;
  RECT 0.000 9.625 4.600 9.935 ;
  RECT 0.000 11.415 4.600 11.725 ;
  RECT 0.000 13.465 4.600 13.775 ;
  RECT 0.000 15.700 4.600 16.010 ;
  RECT 0.000 17.845 4.600 18.345 ;
  RECT 0.000 21.590 4.600 21.900 ;
  RECT 0.000 22.535 4.600 22.845 ;
  RECT 0.000 23.700 4.600 24.010 ;
  RECT 0.000 25.860 4.600 26.230 ;
  RECT 293.805 159.195 298.405 159.265 ;
  RECT 293.805 159.635 298.405 159.775 ;
  RECT 293.805 158.195 298.405 158.255 ;
  RECT 293.805 159.135 298.405 159.195 ;
  RECT 293.805 158.635 298.405 158.755 ;
  RECT 293.805 157.195 298.405 157.255 ;
  RECT 293.805 158.135 298.405 158.195 ;
  RECT 293.805 157.635 298.405 157.755 ;
  RECT 293.805 156.195 298.405 156.255 ;
  RECT 293.805 157.135 298.405 157.195 ;
  RECT 293.805 156.635 298.405 156.755 ;
  RECT 293.805 155.195 298.405 155.255 ;
  RECT 293.805 156.135 298.405 156.195 ;
  RECT 293.805 155.635 298.405 155.755 ;
  RECT 293.805 154.195 298.405 154.255 ;
  RECT 293.805 155.135 298.405 155.195 ;
  RECT 293.805 154.635 298.405 154.755 ;
  RECT 293.805 153.195 298.405 153.255 ;
  RECT 293.805 154.135 298.405 154.195 ;
  RECT 293.805 153.635 298.405 153.755 ;
  RECT 293.805 152.195 298.405 152.255 ;
  RECT 293.805 153.135 298.405 153.195 ;
  RECT 293.805 152.635 298.405 152.755 ;
  RECT 293.805 151.195 298.405 151.255 ;
  RECT 293.805 152.135 298.405 152.195 ;
  RECT 293.805 151.635 298.405 151.755 ;
  RECT 293.805 150.195 298.405 150.255 ;
  RECT 293.805 151.135 298.405 151.195 ;
  RECT 293.805 150.635 298.405 150.755 ;
  RECT 293.805 149.195 298.405 149.255 ;
  RECT 293.805 150.135 298.405 150.195 ;
  RECT 293.805 149.635 298.405 149.755 ;
  RECT 293.805 148.195 298.405 148.255 ;
  RECT 293.805 149.135 298.405 149.195 ;
  RECT 293.805 148.635 298.405 148.755 ;
  RECT 293.805 147.195 298.405 147.255 ;
  RECT 293.805 148.135 298.405 148.195 ;
  RECT 293.805 147.635 298.405 147.755 ;
  RECT 293.805 146.195 298.405 146.255 ;
  RECT 293.805 147.135 298.405 147.195 ;
  RECT 293.805 146.635 298.405 146.755 ;
  RECT 293.805 145.195 298.405 145.255 ;
  RECT 293.805 146.135 298.405 146.195 ;
  RECT 293.805 145.635 298.405 145.755 ;
  RECT 293.805 144.195 298.405 144.255 ;
  RECT 293.805 145.135 298.405 145.195 ;
  RECT 293.805 144.635 298.405 144.755 ;
  RECT 293.805 143.195 298.405 143.255 ;
  RECT 293.805 144.135 298.405 144.195 ;
  RECT 293.805 143.635 298.405 143.755 ;
  RECT 293.805 142.195 298.405 142.255 ;
  RECT 293.805 143.135 298.405 143.195 ;
  RECT 293.805 142.635 298.405 142.755 ;
  RECT 293.805 141.195 298.405 141.255 ;
  RECT 293.805 142.135 298.405 142.195 ;
  RECT 293.805 141.635 298.405 141.755 ;
  RECT 293.805 140.195 298.405 140.255 ;
  RECT 293.805 141.135 298.405 141.195 ;
  RECT 293.805 140.635 298.405 140.755 ;
  RECT 293.805 139.195 298.405 139.255 ;
  RECT 293.805 140.135 298.405 140.195 ;
  RECT 293.805 139.635 298.405 139.755 ;
  RECT 293.805 138.195 298.405 138.255 ;
  RECT 293.805 139.135 298.405 139.195 ;
  RECT 293.805 138.635 298.405 138.755 ;
  RECT 293.805 137.195 298.405 137.255 ;
  RECT 293.805 138.135 298.405 138.195 ;
  RECT 293.805 137.635 298.405 137.755 ;
  RECT 293.805 136.195 298.405 136.255 ;
  RECT 293.805 137.135 298.405 137.195 ;
  RECT 293.805 136.635 298.405 136.755 ;
  RECT 293.805 135.195 298.405 135.255 ;
  RECT 293.805 136.135 298.405 136.195 ;
  RECT 293.805 135.635 298.405 135.755 ;
  RECT 293.805 134.195 298.405 134.255 ;
  RECT 293.805 135.135 298.405 135.195 ;
  RECT 293.805 134.635 298.405 134.755 ;
  RECT 293.805 133.195 298.405 133.255 ;
  RECT 293.805 134.135 298.405 134.195 ;
  RECT 293.805 133.635 298.405 133.755 ;
  RECT 293.805 132.195 298.405 132.255 ;
  RECT 293.805 133.135 298.405 133.195 ;
  RECT 293.805 132.635 298.405 132.755 ;
  RECT 293.805 131.195 298.405 131.255 ;
  RECT 293.805 132.135 298.405 132.195 ;
  RECT 293.805 131.635 298.405 131.755 ;
  RECT 293.805 130.195 298.405 130.255 ;
  RECT 293.805 131.135 298.405 131.195 ;
  RECT 293.805 130.635 298.405 130.755 ;
  RECT 293.805 129.195 298.405 129.255 ;
  RECT 293.805 130.135 298.405 130.195 ;
  RECT 293.805 129.635 298.405 129.755 ;
  RECT 293.805 128.195 298.405 128.255 ;
  RECT 293.805 129.135 298.405 129.195 ;
  RECT 293.805 128.635 298.405 128.755 ;
  RECT 293.805 127.195 298.405 127.255 ;
  RECT 293.805 128.135 298.405 128.195 ;
  RECT 293.805 127.635 298.405 127.755 ;
  RECT 293.805 127.125 298.405 127.195 ;
  RECT 293.805 126.395 298.405 126.465 ;
  RECT 293.805 126.595 298.405 126.735 ;
  RECT 293.805 125.395 298.405 125.455 ;
  RECT 293.805 126.335 298.405 126.395 ;
  RECT 293.805 125.835 298.405 125.955 ;
  RECT 293.805 124.395 298.405 124.455 ;
  RECT 293.805 125.335 298.405 125.395 ;
  RECT 293.805 124.835 298.405 124.955 ;
  RECT 293.805 123.395 298.405 123.455 ;
  RECT 293.805 124.335 298.405 124.395 ;
  RECT 293.805 123.835 298.405 123.955 ;
  RECT 293.805 122.395 298.405 122.455 ;
  RECT 293.805 123.335 298.405 123.395 ;
  RECT 293.805 122.835 298.405 122.955 ;
  RECT 293.805 121.395 298.405 121.455 ;
  RECT 293.805 122.335 298.405 122.395 ;
  RECT 293.805 121.835 298.405 121.955 ;
  RECT 293.805 120.395 298.405 120.455 ;
  RECT 293.805 121.335 298.405 121.395 ;
  RECT 293.805 120.835 298.405 120.955 ;
  RECT 293.805 119.395 298.405 119.455 ;
  RECT 293.805 120.335 298.405 120.395 ;
  RECT 293.805 119.835 298.405 119.955 ;
  RECT 293.805 118.395 298.405 118.455 ;
  RECT 293.805 119.335 298.405 119.395 ;
  RECT 293.805 118.835 298.405 118.955 ;
  RECT 293.805 117.395 298.405 117.455 ;
  RECT 293.805 118.335 298.405 118.395 ;
  RECT 293.805 117.835 298.405 117.955 ;
  RECT 293.805 116.395 298.405 116.455 ;
  RECT 293.805 117.335 298.405 117.395 ;
  RECT 293.805 116.835 298.405 116.955 ;
  RECT 293.805 115.395 298.405 115.455 ;
  RECT 293.805 116.335 298.405 116.395 ;
  RECT 293.805 115.835 298.405 115.955 ;
  RECT 293.805 114.395 298.405 114.455 ;
  RECT 293.805 115.335 298.405 115.395 ;
  RECT 293.805 114.835 298.405 114.955 ;
  RECT 293.805 113.395 298.405 113.455 ;
  RECT 293.805 114.335 298.405 114.395 ;
  RECT 293.805 113.835 298.405 113.955 ;
  RECT 293.805 112.395 298.405 112.455 ;
  RECT 293.805 113.335 298.405 113.395 ;
  RECT 293.805 112.835 298.405 112.955 ;
  RECT 293.805 111.395 298.405 111.455 ;
  RECT 293.805 112.335 298.405 112.395 ;
  RECT 293.805 111.835 298.405 111.955 ;
  RECT 293.805 110.395 298.405 110.455 ;
  RECT 293.805 111.335 298.405 111.395 ;
  RECT 293.805 110.835 298.405 110.955 ;
  RECT 293.805 109.395 298.405 109.455 ;
  RECT 293.805 110.335 298.405 110.395 ;
  RECT 293.805 109.835 298.405 109.955 ;
  RECT 293.805 108.395 298.405 108.455 ;
  RECT 293.805 109.335 298.405 109.395 ;
  RECT 293.805 108.835 298.405 108.955 ;
  RECT 293.805 107.395 298.405 107.455 ;
  RECT 293.805 108.335 298.405 108.395 ;
  RECT 293.805 107.835 298.405 107.955 ;
  RECT 293.805 106.395 298.405 106.455 ;
  RECT 293.805 107.335 298.405 107.395 ;
  RECT 293.805 106.835 298.405 106.955 ;
  RECT 293.805 105.395 298.405 105.455 ;
  RECT 293.805 106.335 298.405 106.395 ;
  RECT 293.805 105.835 298.405 105.955 ;
  RECT 293.805 104.395 298.405 104.455 ;
  RECT 293.805 105.335 298.405 105.395 ;
  RECT 293.805 104.835 298.405 104.955 ;
  RECT 293.805 103.395 298.405 103.455 ;
  RECT 293.805 104.335 298.405 104.395 ;
  RECT 293.805 103.835 298.405 103.955 ;
  RECT 293.805 102.395 298.405 102.455 ;
  RECT 293.805 103.335 298.405 103.395 ;
  RECT 293.805 102.835 298.405 102.955 ;
  RECT 293.805 101.395 298.405 101.455 ;
  RECT 293.805 102.335 298.405 102.395 ;
  RECT 293.805 101.835 298.405 101.955 ;
  RECT 293.805 100.395 298.405 100.455 ;
  RECT 293.805 101.335 298.405 101.395 ;
  RECT 293.805 100.835 298.405 100.955 ;
  RECT 293.805 99.395 298.405 99.455 ;
  RECT 293.805 100.335 298.405 100.395 ;
  RECT 293.805 99.835 298.405 99.955 ;
  RECT 293.805 98.395 298.405 98.455 ;
  RECT 293.805 99.335 298.405 99.395 ;
  RECT 293.805 98.835 298.405 98.955 ;
  RECT 293.805 97.395 298.405 97.455 ;
  RECT 293.805 98.335 298.405 98.395 ;
  RECT 293.805 97.835 298.405 97.955 ;
  RECT 293.805 96.395 298.405 96.455 ;
  RECT 293.805 97.335 298.405 97.395 ;
  RECT 293.805 96.835 298.405 96.955 ;
  RECT 293.805 95.395 298.405 95.455 ;
  RECT 293.805 96.335 298.405 96.395 ;
  RECT 293.805 95.835 298.405 95.955 ;
  RECT 293.805 94.395 298.405 94.455 ;
  RECT 293.805 95.335 298.405 95.395 ;
  RECT 293.805 94.835 298.405 94.955 ;
  RECT 293.805 94.325 298.405 94.395 ;
  RECT 293.805 93.595 298.405 93.665 ;
  RECT 293.805 93.795 298.405 93.935 ;
  RECT 293.805 92.595 298.405 92.655 ;
  RECT 293.805 93.535 298.405 93.595 ;
  RECT 293.805 93.035 298.405 93.155 ;
  RECT 293.805 91.595 298.405 91.655 ;
  RECT 293.805 92.535 298.405 92.595 ;
  RECT 293.805 92.035 298.405 92.155 ;
  RECT 293.805 90.595 298.405 90.655 ;
  RECT 293.805 91.535 298.405 91.595 ;
  RECT 293.805 91.035 298.405 91.155 ;
  RECT 293.805 89.595 298.405 89.655 ;
  RECT 293.805 90.535 298.405 90.595 ;
  RECT 293.805 90.035 298.405 90.155 ;
  RECT 293.805 88.595 298.405 88.655 ;
  RECT 293.805 89.535 298.405 89.595 ;
  RECT 293.805 89.035 298.405 89.155 ;
  RECT 293.805 87.595 298.405 87.655 ;
  RECT 293.805 88.535 298.405 88.595 ;
  RECT 293.805 88.035 298.405 88.155 ;
  RECT 293.805 86.595 298.405 86.655 ;
  RECT 293.805 87.535 298.405 87.595 ;
  RECT 293.805 87.035 298.405 87.155 ;
  RECT 293.805 85.595 298.405 85.655 ;
  RECT 293.805 86.535 298.405 86.595 ;
  RECT 293.805 86.035 298.405 86.155 ;
  RECT 293.805 84.595 298.405 84.655 ;
  RECT 293.805 85.535 298.405 85.595 ;
  RECT 293.805 85.035 298.405 85.155 ;
  RECT 293.805 83.595 298.405 83.655 ;
  RECT 293.805 84.535 298.405 84.595 ;
  RECT 293.805 84.035 298.405 84.155 ;
  RECT 293.805 82.595 298.405 82.655 ;
  RECT 293.805 83.535 298.405 83.595 ;
  RECT 293.805 83.035 298.405 83.155 ;
  RECT 293.805 81.595 298.405 81.655 ;
  RECT 293.805 82.535 298.405 82.595 ;
  RECT 293.805 82.035 298.405 82.155 ;
  RECT 293.805 80.595 298.405 80.655 ;
  RECT 293.805 81.535 298.405 81.595 ;
  RECT 293.805 81.035 298.405 81.155 ;
  RECT 293.805 79.595 298.405 79.655 ;
  RECT 293.805 80.535 298.405 80.595 ;
  RECT 293.805 80.035 298.405 80.155 ;
  RECT 293.805 78.595 298.405 78.655 ;
  RECT 293.805 79.535 298.405 79.595 ;
  RECT 293.805 79.035 298.405 79.155 ;
  RECT 293.805 77.595 298.405 77.655 ;
  RECT 293.805 78.535 298.405 78.595 ;
  RECT 293.805 78.035 298.405 78.155 ;
  RECT 293.805 76.595 298.405 76.655 ;
  RECT 293.805 77.535 298.405 77.595 ;
  RECT 293.805 77.035 298.405 77.155 ;
  RECT 293.805 75.595 298.405 75.655 ;
  RECT 293.805 76.535 298.405 76.595 ;
  RECT 293.805 76.035 298.405 76.155 ;
  RECT 293.805 74.595 298.405 74.655 ;
  RECT 293.805 75.535 298.405 75.595 ;
  RECT 293.805 75.035 298.405 75.155 ;
  RECT 293.805 73.595 298.405 73.655 ;
  RECT 293.805 74.535 298.405 74.595 ;
  RECT 293.805 74.035 298.405 74.155 ;
  RECT 293.805 72.595 298.405 72.655 ;
  RECT 293.805 73.535 298.405 73.595 ;
  RECT 293.805 73.035 298.405 73.155 ;
  RECT 293.805 71.595 298.405 71.655 ;
  RECT 293.805 72.535 298.405 72.595 ;
  RECT 293.805 72.035 298.405 72.155 ;
  RECT 293.805 70.595 298.405 70.655 ;
  RECT 293.805 71.535 298.405 71.595 ;
  RECT 293.805 71.035 298.405 71.155 ;
  RECT 293.805 69.595 298.405 69.655 ;
  RECT 293.805 70.535 298.405 70.595 ;
  RECT 293.805 70.035 298.405 70.155 ;
  RECT 293.805 68.595 298.405 68.655 ;
  RECT 293.805 69.535 298.405 69.595 ;
  RECT 293.805 69.035 298.405 69.155 ;
  RECT 293.805 67.595 298.405 67.655 ;
  RECT 293.805 68.535 298.405 68.595 ;
  RECT 293.805 68.035 298.405 68.155 ;
  RECT 293.805 66.595 298.405 66.655 ;
  RECT 293.805 67.535 298.405 67.595 ;
  RECT 293.805 67.035 298.405 67.155 ;
  RECT 293.805 65.595 298.405 65.655 ;
  RECT 293.805 66.535 298.405 66.595 ;
  RECT 293.805 66.035 298.405 66.155 ;
  RECT 293.805 64.595 298.405 64.655 ;
  RECT 293.805 65.535 298.405 65.595 ;
  RECT 293.805 65.035 298.405 65.155 ;
  RECT 293.805 63.595 298.405 63.655 ;
  RECT 293.805 64.535 298.405 64.595 ;
  RECT 293.805 64.035 298.405 64.155 ;
  RECT 293.805 62.595 298.405 62.655 ;
  RECT 293.805 63.535 298.405 63.595 ;
  RECT 293.805 63.035 298.405 63.155 ;
  RECT 293.805 61.595 298.405 61.655 ;
  RECT 293.805 62.535 298.405 62.595 ;
  RECT 293.805 62.035 298.405 62.155 ;
  RECT 293.805 61.525 298.405 61.595 ;
  RECT 293.805 60.795 298.405 60.865 ;
  RECT 293.805 60.995 298.405 61.135 ;
  RECT 293.805 59.795 298.405 59.855 ;
  RECT 293.805 60.735 298.405 60.795 ;
  RECT 293.805 60.235 298.405 60.355 ;
  RECT 293.805 58.795 298.405 58.855 ;
  RECT 293.805 59.735 298.405 59.795 ;
  RECT 293.805 59.235 298.405 59.355 ;
  RECT 293.805 57.795 298.405 57.855 ;
  RECT 293.805 58.735 298.405 58.795 ;
  RECT 293.805 58.235 298.405 58.355 ;
  RECT 293.805 56.795 298.405 56.855 ;
  RECT 293.805 57.735 298.405 57.795 ;
  RECT 293.805 57.235 298.405 57.355 ;
  RECT 293.805 55.795 298.405 55.855 ;
  RECT 293.805 56.735 298.405 56.795 ;
  RECT 293.805 56.235 298.405 56.355 ;
  RECT 293.805 54.795 298.405 54.855 ;
  RECT 293.805 55.735 298.405 55.795 ;
  RECT 293.805 55.235 298.405 55.355 ;
  RECT 293.805 53.795 298.405 53.855 ;
  RECT 293.805 54.735 298.405 54.795 ;
  RECT 293.805 54.235 298.405 54.355 ;
  RECT 293.805 52.795 298.405 52.855 ;
  RECT 293.805 53.735 298.405 53.795 ;
  RECT 293.805 53.235 298.405 53.355 ;
  RECT 293.805 51.795 298.405 51.855 ;
  RECT 293.805 52.735 298.405 52.795 ;
  RECT 293.805 52.235 298.405 52.355 ;
  RECT 293.805 50.795 298.405 50.855 ;
  RECT 293.805 51.735 298.405 51.795 ;
  RECT 293.805 51.235 298.405 51.355 ;
  RECT 293.805 49.795 298.405 49.855 ;
  RECT 293.805 50.735 298.405 50.795 ;
  RECT 293.805 50.235 298.405 50.355 ;
  RECT 293.805 48.795 298.405 48.855 ;
  RECT 293.805 49.735 298.405 49.795 ;
  RECT 293.805 49.235 298.405 49.355 ;
  RECT 293.805 47.795 298.405 47.855 ;
  RECT 293.805 48.735 298.405 48.795 ;
  RECT 293.805 48.235 298.405 48.355 ;
  RECT 293.805 46.795 298.405 46.855 ;
  RECT 293.805 47.735 298.405 47.795 ;
  RECT 293.805 47.235 298.405 47.355 ;
  RECT 293.805 45.795 298.405 45.855 ;
  RECT 293.805 46.735 298.405 46.795 ;
  RECT 293.805 46.235 298.405 46.355 ;
  RECT 293.805 44.795 298.405 44.855 ;
  RECT 293.805 45.735 298.405 45.795 ;
  RECT 293.805 45.235 298.405 45.355 ;
  RECT 293.805 43.795 298.405 43.855 ;
  RECT 293.805 44.735 298.405 44.795 ;
  RECT 293.805 44.235 298.405 44.355 ;
  RECT 293.805 42.795 298.405 42.855 ;
  RECT 293.805 43.735 298.405 43.795 ;
  RECT 293.805 43.235 298.405 43.355 ;
  RECT 293.805 41.795 298.405 41.855 ;
  RECT 293.805 42.735 298.405 42.795 ;
  RECT 293.805 42.235 298.405 42.355 ;
  RECT 293.805 40.795 298.405 40.855 ;
  RECT 293.805 41.735 298.405 41.795 ;
  RECT 293.805 41.235 298.405 41.355 ;
  RECT 293.805 39.795 298.405 39.855 ;
  RECT 293.805 40.735 298.405 40.795 ;
  RECT 293.805 40.235 298.405 40.355 ;
  RECT 293.805 38.795 298.405 38.855 ;
  RECT 293.805 39.735 298.405 39.795 ;
  RECT 293.805 39.235 298.405 39.355 ;
  RECT 293.805 37.795 298.405 37.855 ;
  RECT 293.805 38.735 298.405 38.795 ;
  RECT 293.805 38.235 298.405 38.355 ;
  RECT 293.805 36.795 298.405 36.855 ;
  RECT 293.805 37.735 298.405 37.795 ;
  RECT 293.805 37.235 298.405 37.355 ;
  RECT 293.805 35.795 298.405 35.855 ;
  RECT 293.805 36.735 298.405 36.795 ;
  RECT 293.805 36.235 298.405 36.355 ;
  RECT 293.805 34.795 298.405 34.855 ;
  RECT 293.805 35.735 298.405 35.795 ;
  RECT 293.805 35.235 298.405 35.355 ;
  RECT 293.805 33.795 298.405 33.855 ;
  RECT 293.805 34.735 298.405 34.795 ;
  RECT 293.805 34.235 298.405 34.355 ;
  RECT 293.805 32.795 298.405 32.855 ;
  RECT 293.805 33.735 298.405 33.795 ;
  RECT 293.805 33.235 298.405 33.355 ;
  RECT 293.805 31.795 298.405 31.855 ;
  RECT 293.805 32.735 298.405 32.795 ;
  RECT 293.805 32.235 298.405 32.355 ;
  RECT 293.805 30.795 298.405 30.855 ;
  RECT 293.805 31.735 298.405 31.795 ;
  RECT 293.805 31.235 298.405 31.355 ;
  RECT 293.805 29.795 298.405 29.855 ;
  RECT 293.805 30.735 298.405 30.795 ;
  RECT 293.805 30.235 298.405 30.355 ;
  RECT 293.805 28.795 298.405 28.855 ;
  RECT 293.805 29.735 298.405 29.795 ;
  RECT 293.805 29.235 298.405 29.355 ;
  RECT 293.805 28.715 298.405 28.795 ;
  RECT 293.805 28.195 298.405 28.335 ;
  RECT 0.000 159.195 4.600 159.265 ;
  RECT 0.000 159.635 4.600 159.775 ;
  RECT 0.000 158.635 4.600 158.755 ;
  RECT 0.000 158.195 4.600 158.255 ;
  RECT 0.000 159.135 4.600 159.195 ;
  RECT 0.000 157.635 4.600 157.755 ;
  RECT 0.000 157.195 4.600 157.255 ;
  RECT 0.000 158.135 4.600 158.195 ;
  RECT 0.000 156.635 4.600 156.755 ;
  RECT 0.000 156.195 4.600 156.255 ;
  RECT 0.000 157.135 4.600 157.195 ;
  RECT 0.000 155.635 4.600 155.755 ;
  RECT 0.000 155.195 4.600 155.255 ;
  RECT 0.000 156.135 4.600 156.195 ;
  RECT 0.000 154.635 4.600 154.755 ;
  RECT 0.000 154.195 4.600 154.255 ;
  RECT 0.000 155.135 4.600 155.195 ;
  RECT 0.000 153.635 4.600 153.755 ;
  RECT 0.000 153.195 4.600 153.255 ;
  RECT 0.000 154.135 4.600 154.195 ;
  RECT 0.000 152.635 4.600 152.755 ;
  RECT 0.000 152.195 4.600 152.255 ;
  RECT 0.000 153.135 4.600 153.195 ;
  RECT 0.000 151.635 4.600 151.755 ;
  RECT 0.000 151.195 4.600 151.255 ;
  RECT 0.000 152.135 4.600 152.195 ;
  RECT 0.000 150.635 4.600 150.755 ;
  RECT 0.000 150.195 4.600 150.255 ;
  RECT 0.000 151.135 4.600 151.195 ;
  RECT 0.000 149.635 4.600 149.755 ;
  RECT 0.000 149.195 4.600 149.255 ;
  RECT 0.000 150.135 4.600 150.195 ;
  RECT 0.000 148.635 4.600 148.755 ;
  RECT 0.000 148.195 4.600 148.255 ;
  RECT 0.000 149.135 4.600 149.195 ;
  RECT 0.000 147.635 4.600 147.755 ;
  RECT 0.000 147.195 4.600 147.255 ;
  RECT 0.000 148.135 4.600 148.195 ;
  RECT 0.000 146.635 4.600 146.755 ;
  RECT 0.000 146.195 4.600 146.255 ;
  RECT 0.000 147.135 4.600 147.195 ;
  RECT 0.000 145.635 4.600 145.755 ;
  RECT 0.000 145.195 4.600 145.255 ;
  RECT 0.000 146.135 4.600 146.195 ;
  RECT 0.000 144.635 4.600 144.755 ;
  RECT 0.000 144.195 4.600 144.255 ;
  RECT 0.000 145.135 4.600 145.195 ;
  RECT 0.000 143.635 4.600 143.755 ;
  RECT 0.000 143.195 4.600 143.255 ;
  RECT 0.000 144.135 4.600 144.195 ;
  RECT 0.000 142.635 4.600 142.755 ;
  RECT 0.000 142.195 4.600 142.255 ;
  RECT 0.000 143.135 4.600 143.195 ;
  RECT 0.000 141.635 4.600 141.755 ;
  RECT 0.000 141.195 4.600 141.255 ;
  RECT 0.000 142.135 4.600 142.195 ;
  RECT 0.000 140.635 4.600 140.755 ;
  RECT 0.000 140.195 4.600 140.255 ;
  RECT 0.000 141.135 4.600 141.195 ;
  RECT 0.000 139.635 4.600 139.755 ;
  RECT 0.000 139.195 4.600 139.255 ;
  RECT 0.000 140.135 4.600 140.195 ;
  RECT 0.000 138.635 4.600 138.755 ;
  RECT 0.000 138.195 4.600 138.255 ;
  RECT 0.000 139.135 4.600 139.195 ;
  RECT 0.000 137.635 4.600 137.755 ;
  RECT 0.000 137.195 4.600 137.255 ;
  RECT 0.000 138.135 4.600 138.195 ;
  RECT 0.000 136.635 4.600 136.755 ;
  RECT 0.000 136.195 4.600 136.255 ;
  RECT 0.000 137.135 4.600 137.195 ;
  RECT 0.000 135.635 4.600 135.755 ;
  RECT 0.000 135.195 4.600 135.255 ;
  RECT 0.000 136.135 4.600 136.195 ;
  RECT 0.000 134.635 4.600 134.755 ;
  RECT 0.000 134.195 4.600 134.255 ;
  RECT 0.000 135.135 4.600 135.195 ;
  RECT 0.000 133.635 4.600 133.755 ;
  RECT 0.000 133.195 4.600 133.255 ;
  RECT 0.000 134.135 4.600 134.195 ;
  RECT 0.000 132.635 4.600 132.755 ;
  RECT 0.000 132.195 4.600 132.255 ;
  RECT 0.000 133.135 4.600 133.195 ;
  RECT 0.000 131.635 4.600 131.755 ;
  RECT 0.000 131.195 4.600 131.255 ;
  RECT 0.000 132.135 4.600 132.195 ;
  RECT 0.000 130.635 4.600 130.755 ;
  RECT 0.000 130.195 4.600 130.255 ;
  RECT 0.000 131.135 4.600 131.195 ;
  RECT 0.000 129.635 4.600 129.755 ;
  RECT 0.000 129.195 4.600 129.255 ;
  RECT 0.000 130.135 4.600 130.195 ;
  RECT 0.000 128.635 4.600 128.755 ;
  RECT 0.000 128.195 4.600 128.255 ;
  RECT 0.000 129.135 4.600 129.195 ;
  RECT 0.000 127.635 4.600 127.755 ;
  RECT 0.000 127.195 4.600 127.255 ;
  RECT 0.000 128.135 4.600 128.195 ;
  RECT 0.000 127.125 4.600 127.195 ;
  RECT 0.000 126.395 4.600 126.465 ;
  RECT 0.000 126.595 4.600 126.735 ;
  RECT 0.000 125.835 4.600 125.955 ;
  RECT 0.000 125.395 4.600 125.455 ;
  RECT 0.000 126.335 4.600 126.395 ;
  RECT 0.000 124.835 4.600 124.955 ;
  RECT 0.000 124.395 4.600 124.455 ;
  RECT 0.000 125.335 4.600 125.395 ;
  RECT 0.000 123.835 4.600 123.955 ;
  RECT 0.000 123.395 4.600 123.455 ;
  RECT 0.000 124.335 4.600 124.395 ;
  RECT 0.000 122.835 4.600 122.955 ;
  RECT 0.000 122.395 4.600 122.455 ;
  RECT 0.000 123.335 4.600 123.395 ;
  RECT 0.000 121.835 4.600 121.955 ;
  RECT 0.000 121.395 4.600 121.455 ;
  RECT 0.000 122.335 4.600 122.395 ;
  RECT 0.000 120.835 4.600 120.955 ;
  RECT 0.000 120.395 4.600 120.455 ;
  RECT 0.000 121.335 4.600 121.395 ;
  RECT 0.000 119.835 4.600 119.955 ;
  RECT 0.000 119.395 4.600 119.455 ;
  RECT 0.000 120.335 4.600 120.395 ;
  RECT 0.000 118.835 4.600 118.955 ;
  RECT 0.000 118.395 4.600 118.455 ;
  RECT 0.000 119.335 4.600 119.395 ;
  RECT 0.000 117.835 4.600 117.955 ;
  RECT 0.000 117.395 4.600 117.455 ;
  RECT 0.000 118.335 4.600 118.395 ;
  RECT 0.000 116.835 4.600 116.955 ;
  RECT 0.000 116.395 4.600 116.455 ;
  RECT 0.000 117.335 4.600 117.395 ;
  RECT 0.000 115.835 4.600 115.955 ;
  RECT 0.000 115.395 4.600 115.455 ;
  RECT 0.000 116.335 4.600 116.395 ;
  RECT 0.000 114.835 4.600 114.955 ;
  RECT 0.000 114.395 4.600 114.455 ;
  RECT 0.000 115.335 4.600 115.395 ;
  RECT 0.000 113.835 4.600 113.955 ;
  RECT 0.000 113.395 4.600 113.455 ;
  RECT 0.000 114.335 4.600 114.395 ;
  RECT 0.000 112.835 4.600 112.955 ;
  RECT 0.000 112.395 4.600 112.455 ;
  RECT 0.000 113.335 4.600 113.395 ;
  RECT 0.000 111.835 4.600 111.955 ;
  RECT 0.000 111.395 4.600 111.455 ;
  RECT 0.000 112.335 4.600 112.395 ;
  RECT 0.000 110.835 4.600 110.955 ;
  RECT 0.000 110.395 4.600 110.455 ;
  RECT 0.000 111.335 4.600 111.395 ;
  RECT 0.000 109.835 4.600 109.955 ;
  RECT 0.000 109.395 4.600 109.455 ;
  RECT 0.000 110.335 4.600 110.395 ;
  RECT 0.000 108.835 4.600 108.955 ;
  RECT 0.000 108.395 4.600 108.455 ;
  RECT 0.000 109.335 4.600 109.395 ;
  RECT 0.000 107.835 4.600 107.955 ;
  RECT 0.000 107.395 4.600 107.455 ;
  RECT 0.000 108.335 4.600 108.395 ;
  RECT 0.000 106.835 4.600 106.955 ;
  RECT 0.000 106.395 4.600 106.455 ;
  RECT 0.000 107.335 4.600 107.395 ;
  RECT 0.000 105.835 4.600 105.955 ;
  RECT 0.000 105.395 4.600 105.455 ;
  RECT 0.000 106.335 4.600 106.395 ;
  RECT 0.000 104.835 4.600 104.955 ;
  RECT 0.000 104.395 4.600 104.455 ;
  RECT 0.000 105.335 4.600 105.395 ;
  RECT 0.000 103.835 4.600 103.955 ;
  RECT 0.000 103.395 4.600 103.455 ;
  RECT 0.000 104.335 4.600 104.395 ;
  RECT 0.000 102.835 4.600 102.955 ;
  RECT 0.000 102.395 4.600 102.455 ;
  RECT 0.000 103.335 4.600 103.395 ;
  RECT 0.000 101.835 4.600 101.955 ;
  RECT 0.000 101.395 4.600 101.455 ;
  RECT 0.000 102.335 4.600 102.395 ;
  RECT 0.000 100.835 4.600 100.955 ;
  RECT 0.000 100.395 4.600 100.455 ;
  RECT 0.000 101.335 4.600 101.395 ;
  RECT 0.000 99.835 4.600 99.955 ;
  RECT 0.000 99.395 4.600 99.455 ;
  RECT 0.000 100.335 4.600 100.395 ;
  RECT 0.000 98.835 4.600 98.955 ;
  RECT 0.000 98.395 4.600 98.455 ;
  RECT 0.000 99.335 4.600 99.395 ;
  RECT 0.000 97.835 4.600 97.955 ;
  RECT 0.000 97.395 4.600 97.455 ;
  RECT 0.000 98.335 4.600 98.395 ;
  RECT 0.000 96.835 4.600 96.955 ;
  RECT 0.000 96.395 4.600 96.455 ;
  RECT 0.000 97.335 4.600 97.395 ;
  RECT 0.000 95.835 4.600 95.955 ;
  RECT 0.000 95.395 4.600 95.455 ;
  RECT 0.000 96.335 4.600 96.395 ;
  RECT 0.000 94.835 4.600 94.955 ;
  RECT 0.000 94.395 4.600 94.455 ;
  RECT 0.000 95.335 4.600 95.395 ;
  RECT 0.000 94.325 4.600 94.395 ;
  RECT 0.000 93.595 4.600 93.665 ;
  RECT 0.000 93.795 4.600 93.935 ;
  RECT 0.000 93.035 4.600 93.155 ;
  RECT 0.000 92.595 4.600 92.655 ;
  RECT 0.000 93.535 4.600 93.595 ;
  RECT 0.000 92.035 4.600 92.155 ;
  RECT 0.000 91.595 4.600 91.655 ;
  RECT 0.000 92.535 4.600 92.595 ;
  RECT 0.000 91.035 4.600 91.155 ;
  RECT 0.000 90.595 4.600 90.655 ;
  RECT 0.000 91.535 4.600 91.595 ;
  RECT 0.000 90.035 4.600 90.155 ;
  RECT 0.000 89.595 4.600 89.655 ;
  RECT 0.000 90.535 4.600 90.595 ;
  RECT 0.000 89.035 4.600 89.155 ;
  RECT 0.000 88.595 4.600 88.655 ;
  RECT 0.000 89.535 4.600 89.595 ;
  RECT 0.000 88.035 4.600 88.155 ;
  RECT 0.000 87.595 4.600 87.655 ;
  RECT 0.000 88.535 4.600 88.595 ;
  RECT 0.000 87.035 4.600 87.155 ;
  RECT 0.000 86.595 4.600 86.655 ;
  RECT 0.000 87.535 4.600 87.595 ;
  RECT 0.000 86.035 4.600 86.155 ;
  RECT 0.000 85.595 4.600 85.655 ;
  RECT 0.000 86.535 4.600 86.595 ;
  RECT 0.000 85.035 4.600 85.155 ;
  RECT 0.000 84.595 4.600 84.655 ;
  RECT 0.000 85.535 4.600 85.595 ;
  RECT 0.000 84.035 4.600 84.155 ;
  RECT 0.000 83.595 4.600 83.655 ;
  RECT 0.000 84.535 4.600 84.595 ;
  RECT 0.000 83.035 4.600 83.155 ;
  RECT 0.000 82.595 4.600 82.655 ;
  RECT 0.000 83.535 4.600 83.595 ;
  RECT 0.000 82.035 4.600 82.155 ;
  RECT 0.000 81.595 4.600 81.655 ;
  RECT 0.000 82.535 4.600 82.595 ;
  RECT 0.000 81.035 4.600 81.155 ;
  RECT 0.000 80.595 4.600 80.655 ;
  RECT 0.000 81.535 4.600 81.595 ;
  RECT 0.000 80.035 4.600 80.155 ;
  RECT 0.000 79.595 4.600 79.655 ;
  RECT 0.000 80.535 4.600 80.595 ;
  RECT 0.000 79.035 4.600 79.155 ;
  RECT 0.000 78.595 4.600 78.655 ;
  RECT 0.000 79.535 4.600 79.595 ;
  RECT 0.000 78.035 4.600 78.155 ;
  RECT 0.000 77.595 4.600 77.655 ;
  RECT 0.000 78.535 4.600 78.595 ;
  RECT 0.000 77.035 4.600 77.155 ;
  RECT 0.000 76.595 4.600 76.655 ;
  RECT 0.000 77.535 4.600 77.595 ;
  RECT 0.000 76.035 4.600 76.155 ;
  RECT 0.000 75.595 4.600 75.655 ;
  RECT 0.000 76.535 4.600 76.595 ;
  RECT 0.000 75.035 4.600 75.155 ;
  RECT 0.000 74.595 4.600 74.655 ;
  RECT 0.000 75.535 4.600 75.595 ;
  RECT 0.000 74.035 4.600 74.155 ;
  RECT 0.000 73.595 4.600 73.655 ;
  RECT 0.000 74.535 4.600 74.595 ;
  RECT 0.000 73.035 4.600 73.155 ;
  RECT 0.000 72.595 4.600 72.655 ;
  RECT 0.000 73.535 4.600 73.595 ;
  RECT 0.000 72.035 4.600 72.155 ;
  RECT 0.000 71.595 4.600 71.655 ;
  RECT 0.000 72.535 4.600 72.595 ;
  RECT 0.000 71.035 4.600 71.155 ;
  RECT 0.000 70.595 4.600 70.655 ;
  RECT 0.000 71.535 4.600 71.595 ;
  RECT 0.000 70.035 4.600 70.155 ;
  RECT 0.000 69.595 4.600 69.655 ;
  RECT 0.000 70.535 4.600 70.595 ;
  RECT 0.000 69.035 4.600 69.155 ;
  RECT 0.000 68.595 4.600 68.655 ;
  RECT 0.000 69.535 4.600 69.595 ;
  RECT 0.000 68.035 4.600 68.155 ;
  RECT 0.000 67.595 4.600 67.655 ;
  RECT 0.000 68.535 4.600 68.595 ;
  RECT 0.000 67.035 4.600 67.155 ;
  RECT 0.000 66.595 4.600 66.655 ;
  RECT 0.000 67.535 4.600 67.595 ;
  RECT 0.000 66.035 4.600 66.155 ;
  RECT 0.000 65.595 4.600 65.655 ;
  RECT 0.000 66.535 4.600 66.595 ;
  RECT 0.000 65.035 4.600 65.155 ;
  RECT 0.000 64.595 4.600 64.655 ;
  RECT 0.000 65.535 4.600 65.595 ;
  RECT 0.000 64.035 4.600 64.155 ;
  RECT 0.000 63.595 4.600 63.655 ;
  RECT 0.000 64.535 4.600 64.595 ;
  RECT 0.000 63.035 4.600 63.155 ;
  RECT 0.000 62.595 4.600 62.655 ;
  RECT 0.000 63.535 4.600 63.595 ;
  RECT 0.000 62.035 4.600 62.155 ;
  RECT 0.000 61.595 4.600 61.655 ;
  RECT 0.000 62.535 4.600 62.595 ;
  RECT 0.000 61.525 4.600 61.595 ;
  RECT 0.000 60.795 4.600 60.865 ;
  RECT 0.000 60.995 4.600 61.135 ;
  RECT 0.000 60.235 4.600 60.355 ;
  RECT 0.000 59.795 4.600 59.855 ;
  RECT 0.000 60.735 4.600 60.795 ;
  RECT 0.000 59.235 4.600 59.355 ;
  RECT 0.000 58.795 4.600 58.855 ;
  RECT 0.000 59.735 4.600 59.795 ;
  RECT 0.000 58.235 4.600 58.355 ;
  RECT 0.000 57.795 4.600 57.855 ;
  RECT 0.000 58.735 4.600 58.795 ;
  RECT 0.000 57.235 4.600 57.355 ;
  RECT 0.000 56.795 4.600 56.855 ;
  RECT 0.000 57.735 4.600 57.795 ;
  RECT 0.000 56.235 4.600 56.355 ;
  RECT 0.000 55.795 4.600 55.855 ;
  RECT 0.000 56.735 4.600 56.795 ;
  RECT 0.000 55.235 4.600 55.355 ;
  RECT 0.000 54.795 4.600 54.855 ;
  RECT 0.000 55.735 4.600 55.795 ;
  RECT 0.000 54.235 4.600 54.355 ;
  RECT 0.000 53.795 4.600 53.855 ;
  RECT 0.000 54.735 4.600 54.795 ;
  RECT 0.000 53.235 4.600 53.355 ;
  RECT 0.000 52.795 4.600 52.855 ;
  RECT 0.000 53.735 4.600 53.795 ;
  RECT 0.000 52.235 4.600 52.355 ;
  RECT 0.000 51.795 4.600 51.855 ;
  RECT 0.000 52.735 4.600 52.795 ;
  RECT 0.000 51.235 4.600 51.355 ;
  RECT 0.000 50.795 4.600 50.855 ;
  RECT 0.000 51.735 4.600 51.795 ;
  RECT 0.000 50.235 4.600 50.355 ;
  RECT 0.000 49.795 4.600 49.855 ;
  RECT 0.000 50.735 4.600 50.795 ;
  RECT 0.000 49.235 4.600 49.355 ;
  RECT 0.000 48.795 4.600 48.855 ;
  RECT 0.000 49.735 4.600 49.795 ;
  RECT 0.000 48.235 4.600 48.355 ;
  RECT 0.000 47.795 4.600 47.855 ;
  RECT 0.000 48.735 4.600 48.795 ;
  RECT 0.000 47.235 4.600 47.355 ;
  RECT 0.000 46.795 4.600 46.855 ;
  RECT 0.000 47.735 4.600 47.795 ;
  RECT 0.000 46.235 4.600 46.355 ;
  RECT 0.000 45.795 4.600 45.855 ;
  RECT 0.000 46.735 4.600 46.795 ;
  RECT 0.000 45.235 4.600 45.355 ;
  RECT 0.000 44.795 4.600 44.855 ;
  RECT 0.000 45.735 4.600 45.795 ;
  RECT 0.000 44.235 4.600 44.355 ;
  RECT 0.000 43.795 4.600 43.855 ;
  RECT 0.000 44.735 4.600 44.795 ;
  RECT 0.000 43.235 4.600 43.355 ;
  RECT 0.000 42.795 4.600 42.855 ;
  RECT 0.000 43.735 4.600 43.795 ;
  RECT 0.000 42.235 4.600 42.355 ;
  RECT 0.000 41.795 4.600 41.855 ;
  RECT 0.000 42.735 4.600 42.795 ;
  RECT 0.000 41.235 4.600 41.355 ;
  RECT 0.000 40.795 4.600 40.855 ;
  RECT 0.000 41.735 4.600 41.795 ;
  RECT 0.000 40.235 4.600 40.355 ;
  RECT 0.000 39.795 4.600 39.855 ;
  RECT 0.000 40.735 4.600 40.795 ;
  RECT 0.000 39.235 4.600 39.355 ;
  RECT 0.000 38.795 4.600 38.855 ;
  RECT 0.000 39.735 4.600 39.795 ;
  RECT 0.000 38.235 4.600 38.355 ;
  RECT 0.000 37.795 4.600 37.855 ;
  RECT 0.000 38.735 4.600 38.795 ;
  RECT 0.000 37.235 4.600 37.355 ;
  RECT 0.000 36.795 4.600 36.855 ;
  RECT 0.000 37.735 4.600 37.795 ;
  RECT 0.000 36.235 4.600 36.355 ;
  RECT 0.000 35.795 4.600 35.855 ;
  RECT 0.000 36.735 4.600 36.795 ;
  RECT 0.000 35.235 4.600 35.355 ;
  RECT 0.000 34.795 4.600 34.855 ;
  RECT 0.000 35.735 4.600 35.795 ;
  RECT 0.000 34.235 4.600 34.355 ;
  RECT 0.000 33.795 4.600 33.855 ;
  RECT 0.000 34.735 4.600 34.795 ;
  RECT 0.000 33.235 4.600 33.355 ;
  RECT 0.000 32.795 4.600 32.855 ;
  RECT 0.000 33.735 4.600 33.795 ;
  RECT 0.000 32.235 4.600 32.355 ;
  RECT 0.000 31.795 4.600 31.855 ;
  RECT 0.000 32.735 4.600 32.795 ;
  RECT 0.000 31.235 4.600 31.355 ;
  RECT 0.000 30.795 4.600 30.855 ;
  RECT 0.000 31.735 4.600 31.795 ;
  RECT 0.000 30.235 4.600 30.355 ;
  RECT 0.000 29.795 4.600 29.855 ;
  RECT 0.000 30.735 4.600 30.795 ;
  RECT 0.000 29.235 4.600 29.355 ;
  RECT 0.000 28.795 4.600 28.855 ;
  RECT 0.000 29.735 4.600 29.795 ;
  RECT 0.000 28.715 4.600 28.795 ;
  RECT 0.000 28.195 4.600 28.335 ;
  LAYER ME4 SPACING 0.160 ;
  RECT 4.600 4.600 148.805 160.240 ;
  LAYER ME4 SPACING 0.160 ;
  RECT 148.920 4.600 149.400 160.240 ;
  LAYER ME4 SPACING 0.160 ;
  RECT 151.860 4.600 152.380 160.240 ;
  LAYER ME4 SPACING 0.160 ;
  RECT 152.580 4.600 154.180 160.240 ;
  LAYER ME4 SPACING 0.160 ;
  RECT 154.395 4.600 154.915 160.240 ;
  LAYER ME4 SPACING 0.160 ;
  RECT 156.695 4.600 157.005 160.240 ;
  LAYER ME4 SPACING 0.160 ;
  RECT 157.165 4.600 293.805 160.240 ;
  LAYER VI2 ;
  RECT 159.220 0.000 159.530 2.000 ;
  RECT 158.770 0.000 159.080 2.000 ;
  RECT 160.870 0.000 161.180 2.000 ;
  RECT 161.320 0.000 161.630 2.000 ;
  RECT 162.970 0.000 163.280 2.000 ;
  RECT 163.420 0.000 163.730 2.000 ;
  RECT 165.070 0.000 165.380 2.000 ;
  RECT 165.520 0.000 165.830 2.000 ;
  RECT 167.170 0.000 167.480 2.000 ;
  RECT 167.620 0.000 167.930 2.000 ;
  RECT 169.270 0.000 169.580 2.000 ;
  RECT 169.720 0.000 170.030 2.000 ;
  RECT 171.370 0.000 171.680 2.000 ;
  RECT 171.820 0.000 172.130 2.000 ;
  RECT 173.470 0.000 173.780 2.000 ;
  RECT 173.920 0.000 174.230 2.000 ;
  RECT 175.570 0.000 175.880 2.000 ;
  RECT 176.020 0.000 176.330 2.000 ;
  RECT 177.670 0.000 177.980 2.000 ;
  RECT 178.120 0.000 178.430 2.000 ;
  RECT 179.770 0.000 180.080 2.000 ;
  RECT 180.220 0.000 180.530 2.000 ;
  RECT 181.870 0.000 182.180 2.000 ;
  RECT 182.320 0.000 182.630 2.000 ;
  RECT 183.970 0.000 184.280 2.000 ;
  RECT 184.420 0.000 184.730 2.000 ;
  RECT 186.070 0.000 186.380 2.000 ;
  RECT 186.520 0.000 186.830 2.000 ;
  RECT 188.170 0.000 188.480 2.000 ;
  RECT 188.620 0.000 188.930 2.000 ;
  RECT 190.270 0.000 190.580 2.000 ;
  RECT 190.720 0.000 191.030 2.000 ;
  RECT 192.370 0.000 192.680 2.000 ;
  RECT 192.820 0.000 193.130 2.000 ;
  RECT 194.470 0.000 194.780 2.000 ;
  RECT 194.920 0.000 195.230 2.000 ;
  RECT 196.570 0.000 196.880 2.000 ;
  RECT 197.020 0.000 197.330 2.000 ;
  RECT 198.670 0.000 198.980 2.000 ;
  RECT 199.120 0.000 199.430 2.000 ;
  RECT 200.770 0.000 201.080 2.000 ;
  RECT 201.220 0.000 201.530 2.000 ;
  RECT 202.870 0.000 203.180 2.000 ;
  RECT 203.320 0.000 203.630 2.000 ;
  RECT 204.970 0.000 205.280 2.000 ;
  RECT 205.420 0.000 205.730 2.000 ;
  RECT 207.070 0.000 207.380 2.000 ;
  RECT 207.520 0.000 207.830 2.000 ;
  RECT 209.170 0.000 209.480 2.000 ;
  RECT 209.620 0.000 209.930 2.000 ;
  RECT 211.270 0.000 211.580 2.000 ;
  RECT 211.720 0.000 212.030 2.000 ;
  RECT 213.370 0.000 213.680 2.000 ;
  RECT 213.820 0.000 214.130 2.000 ;
  RECT 215.470 0.000 215.780 2.000 ;
  RECT 215.920 0.000 216.230 2.000 ;
  RECT 217.570 0.000 217.880 2.000 ;
  RECT 218.020 0.000 218.330 2.000 ;
  RECT 219.670 0.000 219.980 2.000 ;
  RECT 220.120 0.000 220.430 2.000 ;
  RECT 221.770 0.000 222.080 2.000 ;
  RECT 222.220 0.000 222.530 2.000 ;
  RECT 223.870 0.000 224.180 2.000 ;
  RECT 224.320 0.000 224.630 2.000 ;
  RECT 226.420 0.000 226.730 2.000 ;
  RECT 225.970 0.000 226.280 2.000 ;
  RECT 228.070 0.000 228.380 2.000 ;
  RECT 228.520 0.000 228.830 2.000 ;
  RECT 230.170 0.000 230.480 2.000 ;
  RECT 230.620 0.000 230.930 2.000 ;
  RECT 232.270 0.000 232.580 2.000 ;
  RECT 232.720 0.000 233.030 2.000 ;
  RECT 234.370 0.000 234.680 2.000 ;
  RECT 234.820 0.000 235.130 2.000 ;
  RECT 236.470 0.000 236.780 2.000 ;
  RECT 236.920 0.000 237.230 2.000 ;
  RECT 238.570 0.000 238.880 2.000 ;
  RECT 239.020 0.000 239.330 2.000 ;
  RECT 240.670 0.000 240.980 2.000 ;
  RECT 241.120 0.000 241.430 2.000 ;
  RECT 242.770 0.000 243.080 2.000 ;
  RECT 243.220 0.000 243.530 2.000 ;
  RECT 244.870 0.000 245.180 2.000 ;
  RECT 245.320 0.000 245.630 2.000 ;
  RECT 246.970 0.000 247.280 2.000 ;
  RECT 247.420 0.000 247.730 2.000 ;
  RECT 249.070 0.000 249.380 2.000 ;
  RECT 249.520 0.000 249.830 2.000 ;
  RECT 251.170 0.000 251.480 2.000 ;
  RECT 251.620 0.000 251.930 2.000 ;
  RECT 253.270 0.000 253.580 2.000 ;
  RECT 253.720 0.000 254.030 2.000 ;
  RECT 255.370 0.000 255.680 2.000 ;
  RECT 255.820 0.000 256.130 2.000 ;
  RECT 257.470 0.000 257.780 2.000 ;
  RECT 257.920 0.000 258.230 2.000 ;
  RECT 259.570 0.000 259.880 2.000 ;
  RECT 260.020 0.000 260.330 2.000 ;
  RECT 261.670 0.000 261.980 2.000 ;
  RECT 262.120 0.000 262.430 2.000 ;
  RECT 263.770 0.000 264.080 2.000 ;
  RECT 264.220 0.000 264.530 2.000 ;
  RECT 265.870 0.000 266.180 2.000 ;
  RECT 266.320 0.000 266.630 2.000 ;
  RECT 267.970 0.000 268.280 2.000 ;
  RECT 268.420 0.000 268.730 2.000 ;
  RECT 270.070 0.000 270.380 2.000 ;
  RECT 270.520 0.000 270.830 2.000 ;
  RECT 272.170 0.000 272.480 2.000 ;
  RECT 272.620 0.000 272.930 2.000 ;
  RECT 274.270 0.000 274.580 2.000 ;
  RECT 274.720 0.000 275.030 2.000 ;
  RECT 276.370 0.000 276.680 2.000 ;
  RECT 276.820 0.000 277.130 2.000 ;
  RECT 278.470 0.000 278.780 2.000 ;
  RECT 278.920 0.000 279.230 2.000 ;
  RECT 280.570 0.000 280.880 2.000 ;
  RECT 281.020 0.000 281.330 2.000 ;
  RECT 282.670 0.000 282.980 2.000 ;
  RECT 283.120 0.000 283.430 2.000 ;
  RECT 284.770 0.000 285.080 2.000 ;
  RECT 285.220 0.000 285.530 2.000 ;
  RECT 286.870 0.000 287.180 2.000 ;
  RECT 287.320 0.000 287.630 2.000 ;
  RECT 288.970 0.000 289.280 2.000 ;
  RECT 289.420 0.000 289.730 2.000 ;
  RECT 291.070 0.000 291.380 2.000 ;
  RECT 291.520 0.000 291.830 2.000 ;
  RECT 292.645 0.000 292.815 2.000 ;
  RECT 157.750 0.000 158.060 2.000 ;
  RECT 152.690 0.000 153.210 2.000 ;
  RECT 148.050 0.000 148.530 2.000 ;
  RECT 146.055 0.000 146.365 2.000 ;
  RECT 145.380 0.000 145.690 2.000 ;
  RECT 143.775 0.000 144.085 2.000 ;
  RECT 143.100 0.000 143.410 2.000 ;
  RECT 141.495 0.000 141.805 2.000 ;
  RECT 140.820 0.000 141.130 2.000 ;
  RECT 5.590 0.000 5.760 2.000 ;
  RECT 6.995 0.000 7.305 2.000 ;
  RECT 6.545 0.000 6.855 2.000 ;
  RECT 8.645 0.000 8.955 2.000 ;
  RECT 9.095 0.000 9.405 2.000 ;
  RECT 10.745 0.000 11.055 2.000 ;
  RECT 11.195 0.000 11.505 2.000 ;
  RECT 12.845 0.000 13.155 2.000 ;
  RECT 13.295 0.000 13.605 2.000 ;
  RECT 14.945 0.000 15.255 2.000 ;
  RECT 15.395 0.000 15.705 2.000 ;
  RECT 17.045 0.000 17.355 2.000 ;
  RECT 17.495 0.000 17.805 2.000 ;
  RECT 19.145 0.000 19.455 2.000 ;
  RECT 19.595 0.000 19.905 2.000 ;
  RECT 21.245 0.000 21.555 2.000 ;
  RECT 21.695 0.000 22.005 2.000 ;
  RECT 23.345 0.000 23.655 2.000 ;
  RECT 23.795 0.000 24.105 2.000 ;
  RECT 25.445 0.000 25.755 2.000 ;
  RECT 25.895 0.000 26.205 2.000 ;
  RECT 27.545 0.000 27.855 2.000 ;
  RECT 27.995 0.000 28.305 2.000 ;
  RECT 29.645 0.000 29.955 2.000 ;
  RECT 30.095 0.000 30.405 2.000 ;
  RECT 31.745 0.000 32.055 2.000 ;
  RECT 32.195 0.000 32.505 2.000 ;
  RECT 33.845 0.000 34.155 2.000 ;
  RECT 34.295 0.000 34.605 2.000 ;
  RECT 35.945 0.000 36.255 2.000 ;
  RECT 36.395 0.000 36.705 2.000 ;
  RECT 38.045 0.000 38.355 2.000 ;
  RECT 38.495 0.000 38.805 2.000 ;
  RECT 40.145 0.000 40.455 2.000 ;
  RECT 40.595 0.000 40.905 2.000 ;
  RECT 42.245 0.000 42.555 2.000 ;
  RECT 42.695 0.000 43.005 2.000 ;
  RECT 44.345 0.000 44.655 2.000 ;
  RECT 44.795 0.000 45.105 2.000 ;
  RECT 46.445 0.000 46.755 2.000 ;
  RECT 46.895 0.000 47.205 2.000 ;
  RECT 48.545 0.000 48.855 2.000 ;
  RECT 48.995 0.000 49.305 2.000 ;
  RECT 50.645 0.000 50.955 2.000 ;
  RECT 51.095 0.000 51.405 2.000 ;
  RECT 52.745 0.000 53.055 2.000 ;
  RECT 53.195 0.000 53.505 2.000 ;
  RECT 54.845 0.000 55.155 2.000 ;
  RECT 55.295 0.000 55.605 2.000 ;
  RECT 56.945 0.000 57.255 2.000 ;
  RECT 57.395 0.000 57.705 2.000 ;
  RECT 59.045 0.000 59.355 2.000 ;
  RECT 59.495 0.000 59.805 2.000 ;
  RECT 61.145 0.000 61.455 2.000 ;
  RECT 61.595 0.000 61.905 2.000 ;
  RECT 63.245 0.000 63.555 2.000 ;
  RECT 63.695 0.000 64.005 2.000 ;
  RECT 65.345 0.000 65.655 2.000 ;
  RECT 65.795 0.000 66.105 2.000 ;
  RECT 67.445 0.000 67.755 2.000 ;
  RECT 67.895 0.000 68.205 2.000 ;
  RECT 69.545 0.000 69.855 2.000 ;
  RECT 69.995 0.000 70.305 2.000 ;
  RECT 71.645 0.000 71.955 2.000 ;
  RECT 72.095 0.000 72.405 2.000 ;
  RECT 74.195 0.000 74.505 2.000 ;
  RECT 73.745 0.000 74.055 2.000 ;
  RECT 75.845 0.000 76.155 2.000 ;
  RECT 76.295 0.000 76.605 2.000 ;
  RECT 77.945 0.000 78.255 2.000 ;
  RECT 78.395 0.000 78.705 2.000 ;
  RECT 80.045 0.000 80.355 2.000 ;
  RECT 80.495 0.000 80.805 2.000 ;
  RECT 82.145 0.000 82.455 2.000 ;
  RECT 82.595 0.000 82.905 2.000 ;
  RECT 84.245 0.000 84.555 2.000 ;
  RECT 84.695 0.000 85.005 2.000 ;
  RECT 86.345 0.000 86.655 2.000 ;
  RECT 86.795 0.000 87.105 2.000 ;
  RECT 88.445 0.000 88.755 2.000 ;
  RECT 88.895 0.000 89.205 2.000 ;
  RECT 90.545 0.000 90.855 2.000 ;
  RECT 90.995 0.000 91.305 2.000 ;
  RECT 92.645 0.000 92.955 2.000 ;
  RECT 93.095 0.000 93.405 2.000 ;
  RECT 94.745 0.000 95.055 2.000 ;
  RECT 95.195 0.000 95.505 2.000 ;
  RECT 96.845 0.000 97.155 2.000 ;
  RECT 97.295 0.000 97.605 2.000 ;
  RECT 98.945 0.000 99.255 2.000 ;
  RECT 99.395 0.000 99.705 2.000 ;
  RECT 101.045 0.000 101.355 2.000 ;
  RECT 101.495 0.000 101.805 2.000 ;
  RECT 103.145 0.000 103.455 2.000 ;
  RECT 103.595 0.000 103.905 2.000 ;
  RECT 105.245 0.000 105.555 2.000 ;
  RECT 105.695 0.000 106.005 2.000 ;
  RECT 107.345 0.000 107.655 2.000 ;
  RECT 107.795 0.000 108.105 2.000 ;
  RECT 109.445 0.000 109.755 2.000 ;
  RECT 109.895 0.000 110.205 2.000 ;
  RECT 111.545 0.000 111.855 2.000 ;
  RECT 111.995 0.000 112.305 2.000 ;
  RECT 113.645 0.000 113.955 2.000 ;
  RECT 114.095 0.000 114.405 2.000 ;
  RECT 115.745 0.000 116.055 2.000 ;
  RECT 116.195 0.000 116.505 2.000 ;
  RECT 117.845 0.000 118.155 2.000 ;
  RECT 118.295 0.000 118.605 2.000 ;
  RECT 119.945 0.000 120.255 2.000 ;
  RECT 120.395 0.000 120.705 2.000 ;
  RECT 122.045 0.000 122.355 2.000 ;
  RECT 122.495 0.000 122.805 2.000 ;
  RECT 124.145 0.000 124.455 2.000 ;
  RECT 124.595 0.000 124.905 2.000 ;
  RECT 126.245 0.000 126.555 2.000 ;
  RECT 126.695 0.000 127.005 2.000 ;
  RECT 128.345 0.000 128.655 2.000 ;
  RECT 128.795 0.000 129.105 2.000 ;
  RECT 130.445 0.000 130.755 2.000 ;
  RECT 130.895 0.000 131.205 2.000 ;
  RECT 132.545 0.000 132.855 2.000 ;
  RECT 132.995 0.000 133.305 2.000 ;
  RECT 134.645 0.000 134.955 2.000 ;
  RECT 135.095 0.000 135.405 2.000 ;
  RECT 136.745 0.000 137.055 2.000 ;
  RECT 137.195 0.000 137.505 2.000 ;
  RECT 138.845 0.000 139.155 2.000 ;
  RECT 139.295 0.000 139.605 2.000 ;
  RECT 157.750 162.840 158.060 164.840 ;
  RECT 292.645 162.840 292.815 164.840 ;
  RECT 156.695 162.840 157.005 164.840 ;
  RECT 155.755 162.840 156.065 164.840 ;
  RECT 152.690 162.840 153.210 164.840 ;
  RECT 151.310 162.840 151.620 164.840 ;
  RECT 150.285 162.840 150.595 164.840 ;
  RECT 149.765 162.840 150.075 164.840 ;
  RECT 148.050 162.840 148.530 164.840 ;
  RECT 143.775 162.840 144.085 164.840 ;
  RECT 143.100 162.840 143.410 164.840 ;
  RECT 141.495 162.840 141.805 164.840 ;
  RECT 140.870 162.840 141.180 164.840 ;
  RECT 146.055 162.840 146.365 164.840 ;
  RECT 145.380 162.840 145.690 164.840 ;
  RECT 5.590 162.840 5.760 164.840 ;
  RECT 296.405 162.840 298.405 164.840 ;
  RECT 296.405 0.000 298.405 2.000 ;
  RECT 0.000 162.840 2.000 164.840 ;
  RECT 0.000 0.000 2.000 2.000 ;
  RECT 294.105 160.540 296.105 162.540 ;
  RECT 294.105 2.300 296.105 4.300 ;
  RECT 2.300 160.540 4.300 162.540 ;
  RECT 2.300 2.300 4.300 4.300 ;
  LAYER VI1 ;
  RECT 296.405 15.700 298.405 16.010 ;
  RECT 296.405 7.030 298.405 7.340 ;
  RECT 296.405 9.625 298.405 9.935 ;
  RECT 296.405 11.415 298.405 11.725 ;
  RECT 296.405 13.465 298.405 13.775 ;
  RECT 296.405 17.845 298.405 18.345 ;
  RECT 296.405 22.535 298.405 22.845 ;
  RECT 296.405 21.590 298.405 21.900 ;
  RECT 296.405 23.700 298.405 24.010 ;
  RECT 296.405 25.860 298.405 26.230 ;
  RECT 0.000 7.030 2.000 7.340 ;
  RECT 0.000 9.625 2.000 9.935 ;
  RECT 0.000 11.415 2.000 11.725 ;
  RECT 0.000 13.465 2.000 13.775 ;
  RECT 0.000 15.700 2.000 16.010 ;
  RECT 0.000 17.845 2.000 18.345 ;
  RECT 0.000 21.590 2.000 21.900 ;
  RECT 0.000 22.535 2.000 22.845 ;
  RECT 0.000 23.700 2.000 24.010 ;
  RECT 0.000 25.860 2.000 26.230 ;
  RECT 296.405 159.195 298.405 159.265 ;
  RECT 296.405 159.635 298.405 159.775 ;
  RECT 296.405 158.195 298.405 158.255 ;
  RECT 296.405 159.135 298.405 159.195 ;
  RECT 296.405 158.635 298.405 158.755 ;
  RECT 296.405 157.195 298.405 157.255 ;
  RECT 296.405 158.135 298.405 158.195 ;
  RECT 296.405 157.635 298.405 157.755 ;
  RECT 296.405 156.195 298.405 156.255 ;
  RECT 296.405 157.135 298.405 157.195 ;
  RECT 296.405 156.635 298.405 156.755 ;
  RECT 296.405 155.195 298.405 155.255 ;
  RECT 296.405 156.135 298.405 156.195 ;
  RECT 296.405 155.635 298.405 155.755 ;
  RECT 296.405 154.195 298.405 154.255 ;
  RECT 296.405 155.135 298.405 155.195 ;
  RECT 296.405 154.635 298.405 154.755 ;
  RECT 296.405 153.195 298.405 153.255 ;
  RECT 296.405 154.135 298.405 154.195 ;
  RECT 296.405 153.635 298.405 153.755 ;
  RECT 296.405 152.195 298.405 152.255 ;
  RECT 296.405 153.135 298.405 153.195 ;
  RECT 296.405 152.635 298.405 152.755 ;
  RECT 296.405 151.195 298.405 151.255 ;
  RECT 296.405 152.135 298.405 152.195 ;
  RECT 296.405 151.635 298.405 151.755 ;
  RECT 296.405 150.195 298.405 150.255 ;
  RECT 296.405 151.135 298.405 151.195 ;
  RECT 296.405 150.635 298.405 150.755 ;
  RECT 296.405 149.195 298.405 149.255 ;
  RECT 296.405 150.135 298.405 150.195 ;
  RECT 296.405 149.635 298.405 149.755 ;
  RECT 296.405 148.195 298.405 148.255 ;
  RECT 296.405 149.135 298.405 149.195 ;
  RECT 296.405 148.635 298.405 148.755 ;
  RECT 296.405 147.195 298.405 147.255 ;
  RECT 296.405 148.135 298.405 148.195 ;
  RECT 296.405 147.635 298.405 147.755 ;
  RECT 296.405 146.195 298.405 146.255 ;
  RECT 296.405 147.135 298.405 147.195 ;
  RECT 296.405 146.635 298.405 146.755 ;
  RECT 296.405 145.195 298.405 145.255 ;
  RECT 296.405 146.135 298.405 146.195 ;
  RECT 296.405 145.635 298.405 145.755 ;
  RECT 296.405 144.195 298.405 144.255 ;
  RECT 296.405 145.135 298.405 145.195 ;
  RECT 296.405 144.635 298.405 144.755 ;
  RECT 296.405 143.195 298.405 143.255 ;
  RECT 296.405 144.135 298.405 144.195 ;
  RECT 296.405 143.635 298.405 143.755 ;
  RECT 296.405 142.195 298.405 142.255 ;
  RECT 296.405 143.135 298.405 143.195 ;
  RECT 296.405 142.635 298.405 142.755 ;
  RECT 296.405 141.195 298.405 141.255 ;
  RECT 296.405 142.135 298.405 142.195 ;
  RECT 296.405 141.635 298.405 141.755 ;
  RECT 296.405 140.195 298.405 140.255 ;
  RECT 296.405 141.135 298.405 141.195 ;
  RECT 296.405 140.635 298.405 140.755 ;
  RECT 296.405 139.195 298.405 139.255 ;
  RECT 296.405 140.135 298.405 140.195 ;
  RECT 296.405 139.635 298.405 139.755 ;
  RECT 296.405 138.195 298.405 138.255 ;
  RECT 296.405 139.135 298.405 139.195 ;
  RECT 296.405 138.635 298.405 138.755 ;
  RECT 296.405 137.195 298.405 137.255 ;
  RECT 296.405 138.135 298.405 138.195 ;
  RECT 296.405 137.635 298.405 137.755 ;
  RECT 296.405 136.195 298.405 136.255 ;
  RECT 296.405 137.135 298.405 137.195 ;
  RECT 296.405 136.635 298.405 136.755 ;
  RECT 296.405 135.195 298.405 135.255 ;
  RECT 296.405 136.135 298.405 136.195 ;
  RECT 296.405 135.635 298.405 135.755 ;
  RECT 296.405 134.195 298.405 134.255 ;
  RECT 296.405 135.135 298.405 135.195 ;
  RECT 296.405 134.635 298.405 134.755 ;
  RECT 296.405 133.195 298.405 133.255 ;
  RECT 296.405 134.135 298.405 134.195 ;
  RECT 296.405 133.635 298.405 133.755 ;
  RECT 296.405 132.195 298.405 132.255 ;
  RECT 296.405 133.135 298.405 133.195 ;
  RECT 296.405 132.635 298.405 132.755 ;
  RECT 296.405 131.195 298.405 131.255 ;
  RECT 296.405 132.135 298.405 132.195 ;
  RECT 296.405 131.635 298.405 131.755 ;
  RECT 296.405 130.195 298.405 130.255 ;
  RECT 296.405 131.135 298.405 131.195 ;
  RECT 296.405 130.635 298.405 130.755 ;
  RECT 296.405 129.195 298.405 129.255 ;
  RECT 296.405 130.135 298.405 130.195 ;
  RECT 296.405 129.635 298.405 129.755 ;
  RECT 296.405 128.195 298.405 128.255 ;
  RECT 296.405 129.135 298.405 129.195 ;
  RECT 296.405 128.635 298.405 128.755 ;
  RECT 296.405 127.195 298.405 127.255 ;
  RECT 296.405 128.135 298.405 128.195 ;
  RECT 296.405 127.635 298.405 127.755 ;
  RECT 296.405 127.125 298.405 127.195 ;
  RECT 296.405 126.395 298.405 126.465 ;
  RECT 296.405 126.595 298.405 126.735 ;
  RECT 296.405 125.395 298.405 125.455 ;
  RECT 296.405 126.335 298.405 126.395 ;
  RECT 296.405 125.835 298.405 125.955 ;
  RECT 296.405 124.395 298.405 124.455 ;
  RECT 296.405 125.335 298.405 125.395 ;
  RECT 296.405 124.835 298.405 124.955 ;
  RECT 296.405 123.395 298.405 123.455 ;
  RECT 296.405 124.335 298.405 124.395 ;
  RECT 296.405 123.835 298.405 123.955 ;
  RECT 296.405 122.395 298.405 122.455 ;
  RECT 296.405 123.335 298.405 123.395 ;
  RECT 296.405 122.835 298.405 122.955 ;
  RECT 296.405 121.395 298.405 121.455 ;
  RECT 296.405 122.335 298.405 122.395 ;
  RECT 296.405 121.835 298.405 121.955 ;
  RECT 296.405 120.395 298.405 120.455 ;
  RECT 296.405 121.335 298.405 121.395 ;
  RECT 296.405 120.835 298.405 120.955 ;
  RECT 296.405 119.395 298.405 119.455 ;
  RECT 296.405 120.335 298.405 120.395 ;
  RECT 296.405 119.835 298.405 119.955 ;
  RECT 296.405 118.395 298.405 118.455 ;
  RECT 296.405 119.335 298.405 119.395 ;
  RECT 296.405 118.835 298.405 118.955 ;
  RECT 296.405 117.395 298.405 117.455 ;
  RECT 296.405 118.335 298.405 118.395 ;
  RECT 296.405 117.835 298.405 117.955 ;
  RECT 296.405 116.395 298.405 116.455 ;
  RECT 296.405 117.335 298.405 117.395 ;
  RECT 296.405 116.835 298.405 116.955 ;
  RECT 296.405 115.395 298.405 115.455 ;
  RECT 296.405 116.335 298.405 116.395 ;
  RECT 296.405 115.835 298.405 115.955 ;
  RECT 296.405 114.395 298.405 114.455 ;
  RECT 296.405 115.335 298.405 115.395 ;
  RECT 296.405 114.835 298.405 114.955 ;
  RECT 296.405 113.395 298.405 113.455 ;
  RECT 296.405 114.335 298.405 114.395 ;
  RECT 296.405 113.835 298.405 113.955 ;
  RECT 296.405 112.395 298.405 112.455 ;
  RECT 296.405 113.335 298.405 113.395 ;
  RECT 296.405 112.835 298.405 112.955 ;
  RECT 296.405 111.395 298.405 111.455 ;
  RECT 296.405 112.335 298.405 112.395 ;
  RECT 296.405 111.835 298.405 111.955 ;
  RECT 296.405 110.395 298.405 110.455 ;
  RECT 296.405 111.335 298.405 111.395 ;
  RECT 296.405 110.835 298.405 110.955 ;
  RECT 296.405 109.395 298.405 109.455 ;
  RECT 296.405 110.335 298.405 110.395 ;
  RECT 296.405 109.835 298.405 109.955 ;
  RECT 296.405 108.395 298.405 108.455 ;
  RECT 296.405 109.335 298.405 109.395 ;
  RECT 296.405 108.835 298.405 108.955 ;
  RECT 296.405 107.395 298.405 107.455 ;
  RECT 296.405 108.335 298.405 108.395 ;
  RECT 296.405 107.835 298.405 107.955 ;
  RECT 296.405 106.395 298.405 106.455 ;
  RECT 296.405 107.335 298.405 107.395 ;
  RECT 296.405 106.835 298.405 106.955 ;
  RECT 296.405 105.395 298.405 105.455 ;
  RECT 296.405 106.335 298.405 106.395 ;
  RECT 296.405 105.835 298.405 105.955 ;
  RECT 296.405 104.395 298.405 104.455 ;
  RECT 296.405 105.335 298.405 105.395 ;
  RECT 296.405 104.835 298.405 104.955 ;
  RECT 296.405 103.395 298.405 103.455 ;
  RECT 296.405 104.335 298.405 104.395 ;
  RECT 296.405 103.835 298.405 103.955 ;
  RECT 296.405 102.395 298.405 102.455 ;
  RECT 296.405 103.335 298.405 103.395 ;
  RECT 296.405 102.835 298.405 102.955 ;
  RECT 296.405 101.395 298.405 101.455 ;
  RECT 296.405 102.335 298.405 102.395 ;
  RECT 296.405 101.835 298.405 101.955 ;
  RECT 296.405 100.395 298.405 100.455 ;
  RECT 296.405 101.335 298.405 101.395 ;
  RECT 296.405 100.835 298.405 100.955 ;
  RECT 296.405 99.395 298.405 99.455 ;
  RECT 296.405 100.335 298.405 100.395 ;
  RECT 296.405 99.835 298.405 99.955 ;
  RECT 296.405 98.395 298.405 98.455 ;
  RECT 296.405 99.335 298.405 99.395 ;
  RECT 296.405 98.835 298.405 98.955 ;
  RECT 296.405 97.395 298.405 97.455 ;
  RECT 296.405 98.335 298.405 98.395 ;
  RECT 296.405 97.835 298.405 97.955 ;
  RECT 296.405 96.395 298.405 96.455 ;
  RECT 296.405 97.335 298.405 97.395 ;
  RECT 296.405 96.835 298.405 96.955 ;
  RECT 296.405 95.395 298.405 95.455 ;
  RECT 296.405 96.335 298.405 96.395 ;
  RECT 296.405 95.835 298.405 95.955 ;
  RECT 296.405 94.395 298.405 94.455 ;
  RECT 296.405 95.335 298.405 95.395 ;
  RECT 296.405 94.835 298.405 94.955 ;
  RECT 296.405 94.325 298.405 94.395 ;
  RECT 296.405 93.595 298.405 93.665 ;
  RECT 296.405 93.795 298.405 93.935 ;
  RECT 296.405 92.595 298.405 92.655 ;
  RECT 296.405 93.535 298.405 93.595 ;
  RECT 296.405 93.035 298.405 93.155 ;
  RECT 296.405 91.595 298.405 91.655 ;
  RECT 296.405 92.535 298.405 92.595 ;
  RECT 296.405 92.035 298.405 92.155 ;
  RECT 296.405 90.595 298.405 90.655 ;
  RECT 296.405 91.535 298.405 91.595 ;
  RECT 296.405 91.035 298.405 91.155 ;
  RECT 296.405 89.595 298.405 89.655 ;
  RECT 296.405 90.535 298.405 90.595 ;
  RECT 296.405 90.035 298.405 90.155 ;
  RECT 296.405 88.595 298.405 88.655 ;
  RECT 296.405 89.535 298.405 89.595 ;
  RECT 296.405 89.035 298.405 89.155 ;
  RECT 296.405 87.595 298.405 87.655 ;
  RECT 296.405 88.535 298.405 88.595 ;
  RECT 296.405 88.035 298.405 88.155 ;
  RECT 296.405 86.595 298.405 86.655 ;
  RECT 296.405 87.535 298.405 87.595 ;
  RECT 296.405 87.035 298.405 87.155 ;
  RECT 296.405 85.595 298.405 85.655 ;
  RECT 296.405 86.535 298.405 86.595 ;
  RECT 296.405 86.035 298.405 86.155 ;
  RECT 296.405 84.595 298.405 84.655 ;
  RECT 296.405 85.535 298.405 85.595 ;
  RECT 296.405 85.035 298.405 85.155 ;
  RECT 296.405 83.595 298.405 83.655 ;
  RECT 296.405 84.535 298.405 84.595 ;
  RECT 296.405 84.035 298.405 84.155 ;
  RECT 296.405 82.595 298.405 82.655 ;
  RECT 296.405 83.535 298.405 83.595 ;
  RECT 296.405 83.035 298.405 83.155 ;
  RECT 296.405 81.595 298.405 81.655 ;
  RECT 296.405 82.535 298.405 82.595 ;
  RECT 296.405 82.035 298.405 82.155 ;
  RECT 296.405 80.595 298.405 80.655 ;
  RECT 296.405 81.535 298.405 81.595 ;
  RECT 296.405 81.035 298.405 81.155 ;
  RECT 296.405 79.595 298.405 79.655 ;
  RECT 296.405 80.535 298.405 80.595 ;
  RECT 296.405 80.035 298.405 80.155 ;
  RECT 296.405 78.595 298.405 78.655 ;
  RECT 296.405 79.535 298.405 79.595 ;
  RECT 296.405 79.035 298.405 79.155 ;
  RECT 296.405 77.595 298.405 77.655 ;
  RECT 296.405 78.535 298.405 78.595 ;
  RECT 296.405 78.035 298.405 78.155 ;
  RECT 296.405 76.595 298.405 76.655 ;
  RECT 296.405 77.535 298.405 77.595 ;
  RECT 296.405 77.035 298.405 77.155 ;
  RECT 296.405 75.595 298.405 75.655 ;
  RECT 296.405 76.535 298.405 76.595 ;
  RECT 296.405 76.035 298.405 76.155 ;
  RECT 296.405 74.595 298.405 74.655 ;
  RECT 296.405 75.535 298.405 75.595 ;
  RECT 296.405 75.035 298.405 75.155 ;
  RECT 296.405 73.595 298.405 73.655 ;
  RECT 296.405 74.535 298.405 74.595 ;
  RECT 296.405 74.035 298.405 74.155 ;
  RECT 296.405 72.595 298.405 72.655 ;
  RECT 296.405 73.535 298.405 73.595 ;
  RECT 296.405 73.035 298.405 73.155 ;
  RECT 296.405 71.595 298.405 71.655 ;
  RECT 296.405 72.535 298.405 72.595 ;
  RECT 296.405 72.035 298.405 72.155 ;
  RECT 296.405 70.595 298.405 70.655 ;
  RECT 296.405 71.535 298.405 71.595 ;
  RECT 296.405 71.035 298.405 71.155 ;
  RECT 296.405 69.595 298.405 69.655 ;
  RECT 296.405 70.535 298.405 70.595 ;
  RECT 296.405 70.035 298.405 70.155 ;
  RECT 296.405 68.595 298.405 68.655 ;
  RECT 296.405 69.535 298.405 69.595 ;
  RECT 296.405 69.035 298.405 69.155 ;
  RECT 296.405 67.595 298.405 67.655 ;
  RECT 296.405 68.535 298.405 68.595 ;
  RECT 296.405 68.035 298.405 68.155 ;
  RECT 296.405 66.595 298.405 66.655 ;
  RECT 296.405 67.535 298.405 67.595 ;
  RECT 296.405 67.035 298.405 67.155 ;
  RECT 296.405 65.595 298.405 65.655 ;
  RECT 296.405 66.535 298.405 66.595 ;
  RECT 296.405 66.035 298.405 66.155 ;
  RECT 296.405 64.595 298.405 64.655 ;
  RECT 296.405 65.535 298.405 65.595 ;
  RECT 296.405 65.035 298.405 65.155 ;
  RECT 296.405 63.595 298.405 63.655 ;
  RECT 296.405 64.535 298.405 64.595 ;
  RECT 296.405 64.035 298.405 64.155 ;
  RECT 296.405 62.595 298.405 62.655 ;
  RECT 296.405 63.535 298.405 63.595 ;
  RECT 296.405 63.035 298.405 63.155 ;
  RECT 296.405 61.595 298.405 61.655 ;
  RECT 296.405 62.535 298.405 62.595 ;
  RECT 296.405 62.035 298.405 62.155 ;
  RECT 296.405 61.525 298.405 61.595 ;
  RECT 296.405 60.795 298.405 60.865 ;
  RECT 296.405 60.995 298.405 61.135 ;
  RECT 296.405 59.795 298.405 59.855 ;
  RECT 296.405 60.735 298.405 60.795 ;
  RECT 296.405 60.235 298.405 60.355 ;
  RECT 296.405 58.795 298.405 58.855 ;
  RECT 296.405 59.735 298.405 59.795 ;
  RECT 296.405 59.235 298.405 59.355 ;
  RECT 296.405 57.795 298.405 57.855 ;
  RECT 296.405 58.735 298.405 58.795 ;
  RECT 296.405 58.235 298.405 58.355 ;
  RECT 296.405 56.795 298.405 56.855 ;
  RECT 296.405 57.735 298.405 57.795 ;
  RECT 296.405 57.235 298.405 57.355 ;
  RECT 296.405 55.795 298.405 55.855 ;
  RECT 296.405 56.735 298.405 56.795 ;
  RECT 296.405 56.235 298.405 56.355 ;
  RECT 296.405 54.795 298.405 54.855 ;
  RECT 296.405 55.735 298.405 55.795 ;
  RECT 296.405 55.235 298.405 55.355 ;
  RECT 296.405 53.795 298.405 53.855 ;
  RECT 296.405 54.735 298.405 54.795 ;
  RECT 296.405 54.235 298.405 54.355 ;
  RECT 296.405 52.795 298.405 52.855 ;
  RECT 296.405 53.735 298.405 53.795 ;
  RECT 296.405 53.235 298.405 53.355 ;
  RECT 296.405 51.795 298.405 51.855 ;
  RECT 296.405 52.735 298.405 52.795 ;
  RECT 296.405 52.235 298.405 52.355 ;
  RECT 296.405 50.795 298.405 50.855 ;
  RECT 296.405 51.735 298.405 51.795 ;
  RECT 296.405 51.235 298.405 51.355 ;
  RECT 296.405 49.795 298.405 49.855 ;
  RECT 296.405 50.735 298.405 50.795 ;
  RECT 296.405 50.235 298.405 50.355 ;
  RECT 296.405 48.795 298.405 48.855 ;
  RECT 296.405 49.735 298.405 49.795 ;
  RECT 296.405 49.235 298.405 49.355 ;
  RECT 296.405 47.795 298.405 47.855 ;
  RECT 296.405 48.735 298.405 48.795 ;
  RECT 296.405 48.235 298.405 48.355 ;
  RECT 296.405 46.795 298.405 46.855 ;
  RECT 296.405 47.735 298.405 47.795 ;
  RECT 296.405 47.235 298.405 47.355 ;
  RECT 296.405 45.795 298.405 45.855 ;
  RECT 296.405 46.735 298.405 46.795 ;
  RECT 296.405 46.235 298.405 46.355 ;
  RECT 296.405 44.795 298.405 44.855 ;
  RECT 296.405 45.735 298.405 45.795 ;
  RECT 296.405 45.235 298.405 45.355 ;
  RECT 296.405 43.795 298.405 43.855 ;
  RECT 296.405 44.735 298.405 44.795 ;
  RECT 296.405 44.235 298.405 44.355 ;
  RECT 296.405 42.795 298.405 42.855 ;
  RECT 296.405 43.735 298.405 43.795 ;
  RECT 296.405 43.235 298.405 43.355 ;
  RECT 296.405 41.795 298.405 41.855 ;
  RECT 296.405 42.735 298.405 42.795 ;
  RECT 296.405 42.235 298.405 42.355 ;
  RECT 296.405 40.795 298.405 40.855 ;
  RECT 296.405 41.735 298.405 41.795 ;
  RECT 296.405 41.235 298.405 41.355 ;
  RECT 296.405 39.795 298.405 39.855 ;
  RECT 296.405 40.735 298.405 40.795 ;
  RECT 296.405 40.235 298.405 40.355 ;
  RECT 296.405 38.795 298.405 38.855 ;
  RECT 296.405 39.735 298.405 39.795 ;
  RECT 296.405 39.235 298.405 39.355 ;
  RECT 296.405 37.795 298.405 37.855 ;
  RECT 296.405 38.735 298.405 38.795 ;
  RECT 296.405 38.235 298.405 38.355 ;
  RECT 296.405 36.795 298.405 36.855 ;
  RECT 296.405 37.735 298.405 37.795 ;
  RECT 296.405 37.235 298.405 37.355 ;
  RECT 296.405 35.795 298.405 35.855 ;
  RECT 296.405 36.735 298.405 36.795 ;
  RECT 296.405 36.235 298.405 36.355 ;
  RECT 296.405 34.795 298.405 34.855 ;
  RECT 296.405 35.735 298.405 35.795 ;
  RECT 296.405 35.235 298.405 35.355 ;
  RECT 296.405 33.795 298.405 33.855 ;
  RECT 296.405 34.735 298.405 34.795 ;
  RECT 296.405 34.235 298.405 34.355 ;
  RECT 296.405 32.795 298.405 32.855 ;
  RECT 296.405 33.735 298.405 33.795 ;
  RECT 296.405 33.235 298.405 33.355 ;
  RECT 296.405 31.795 298.405 31.855 ;
  RECT 296.405 32.735 298.405 32.795 ;
  RECT 296.405 32.235 298.405 32.355 ;
  RECT 296.405 30.795 298.405 30.855 ;
  RECT 296.405 31.735 298.405 31.795 ;
  RECT 296.405 31.235 298.405 31.355 ;
  RECT 296.405 29.795 298.405 29.855 ;
  RECT 296.405 30.735 298.405 30.795 ;
  RECT 296.405 30.235 298.405 30.355 ;
  RECT 296.405 28.795 298.405 28.855 ;
  RECT 296.405 29.735 298.405 29.795 ;
  RECT 296.405 29.235 298.405 29.355 ;
  RECT 296.405 28.715 298.405 28.795 ;
  RECT 296.405 28.195 298.405 28.335 ;
  RECT 0.000 159.195 2.000 159.265 ;
  RECT 0.000 159.635 2.000 159.775 ;
  RECT 0.000 158.635 2.000 158.755 ;
  RECT 0.000 158.195 2.000 158.255 ;
  RECT 0.000 159.135 2.000 159.195 ;
  RECT 0.000 157.635 2.000 157.755 ;
  RECT 0.000 157.195 2.000 157.255 ;
  RECT 0.000 158.135 2.000 158.195 ;
  RECT 0.000 156.635 2.000 156.755 ;
  RECT 0.000 156.195 2.000 156.255 ;
  RECT 0.000 157.135 2.000 157.195 ;
  RECT 0.000 155.635 2.000 155.755 ;
  RECT 0.000 155.195 2.000 155.255 ;
  RECT 0.000 156.135 2.000 156.195 ;
  RECT 0.000 154.635 2.000 154.755 ;
  RECT 0.000 154.195 2.000 154.255 ;
  RECT 0.000 155.135 2.000 155.195 ;
  RECT 0.000 153.635 2.000 153.755 ;
  RECT 0.000 153.195 2.000 153.255 ;
  RECT 0.000 154.135 2.000 154.195 ;
  RECT 0.000 152.635 2.000 152.755 ;
  RECT 0.000 152.195 2.000 152.255 ;
  RECT 0.000 153.135 2.000 153.195 ;
  RECT 0.000 151.635 2.000 151.755 ;
  RECT 0.000 151.195 2.000 151.255 ;
  RECT 0.000 152.135 2.000 152.195 ;
  RECT 0.000 150.635 2.000 150.755 ;
  RECT 0.000 150.195 2.000 150.255 ;
  RECT 0.000 151.135 2.000 151.195 ;
  RECT 0.000 149.635 2.000 149.755 ;
  RECT 0.000 149.195 2.000 149.255 ;
  RECT 0.000 150.135 2.000 150.195 ;
  RECT 0.000 148.635 2.000 148.755 ;
  RECT 0.000 148.195 2.000 148.255 ;
  RECT 0.000 149.135 2.000 149.195 ;
  RECT 0.000 147.635 2.000 147.755 ;
  RECT 0.000 147.195 2.000 147.255 ;
  RECT 0.000 148.135 2.000 148.195 ;
  RECT 0.000 146.635 2.000 146.755 ;
  RECT 0.000 146.195 2.000 146.255 ;
  RECT 0.000 147.135 2.000 147.195 ;
  RECT 0.000 145.635 2.000 145.755 ;
  RECT 0.000 145.195 2.000 145.255 ;
  RECT 0.000 146.135 2.000 146.195 ;
  RECT 0.000 144.635 2.000 144.755 ;
  RECT 0.000 144.195 2.000 144.255 ;
  RECT 0.000 145.135 2.000 145.195 ;
  RECT 0.000 143.635 2.000 143.755 ;
  RECT 0.000 143.195 2.000 143.255 ;
  RECT 0.000 144.135 2.000 144.195 ;
  RECT 0.000 142.635 2.000 142.755 ;
  RECT 0.000 142.195 2.000 142.255 ;
  RECT 0.000 143.135 2.000 143.195 ;
  RECT 0.000 141.635 2.000 141.755 ;
  RECT 0.000 141.195 2.000 141.255 ;
  RECT 0.000 142.135 2.000 142.195 ;
  RECT 0.000 140.635 2.000 140.755 ;
  RECT 0.000 140.195 2.000 140.255 ;
  RECT 0.000 141.135 2.000 141.195 ;
  RECT 0.000 139.635 2.000 139.755 ;
  RECT 0.000 139.195 2.000 139.255 ;
  RECT 0.000 140.135 2.000 140.195 ;
  RECT 0.000 138.635 2.000 138.755 ;
  RECT 0.000 138.195 2.000 138.255 ;
  RECT 0.000 139.135 2.000 139.195 ;
  RECT 0.000 137.635 2.000 137.755 ;
  RECT 0.000 137.195 2.000 137.255 ;
  RECT 0.000 138.135 2.000 138.195 ;
  RECT 0.000 136.635 2.000 136.755 ;
  RECT 0.000 136.195 2.000 136.255 ;
  RECT 0.000 137.135 2.000 137.195 ;
  RECT 0.000 135.635 2.000 135.755 ;
  RECT 0.000 135.195 2.000 135.255 ;
  RECT 0.000 136.135 2.000 136.195 ;
  RECT 0.000 134.635 2.000 134.755 ;
  RECT 0.000 134.195 2.000 134.255 ;
  RECT 0.000 135.135 2.000 135.195 ;
  RECT 0.000 133.635 2.000 133.755 ;
  RECT 0.000 133.195 2.000 133.255 ;
  RECT 0.000 134.135 2.000 134.195 ;
  RECT 0.000 132.635 2.000 132.755 ;
  RECT 0.000 132.195 2.000 132.255 ;
  RECT 0.000 133.135 2.000 133.195 ;
  RECT 0.000 131.635 2.000 131.755 ;
  RECT 0.000 131.195 2.000 131.255 ;
  RECT 0.000 132.135 2.000 132.195 ;
  RECT 0.000 130.635 2.000 130.755 ;
  RECT 0.000 130.195 2.000 130.255 ;
  RECT 0.000 131.135 2.000 131.195 ;
  RECT 0.000 129.635 2.000 129.755 ;
  RECT 0.000 129.195 2.000 129.255 ;
  RECT 0.000 130.135 2.000 130.195 ;
  RECT 0.000 128.635 2.000 128.755 ;
  RECT 0.000 128.195 2.000 128.255 ;
  RECT 0.000 129.135 2.000 129.195 ;
  RECT 0.000 127.635 2.000 127.755 ;
  RECT 0.000 127.195 2.000 127.255 ;
  RECT 0.000 128.135 2.000 128.195 ;
  RECT 0.000 127.125 2.000 127.195 ;
  RECT 0.000 126.395 2.000 126.465 ;
  RECT 0.000 126.595 2.000 126.735 ;
  RECT 0.000 125.835 2.000 125.955 ;
  RECT 0.000 125.395 2.000 125.455 ;
  RECT 0.000 126.335 2.000 126.395 ;
  RECT 0.000 124.835 2.000 124.955 ;
  RECT 0.000 124.395 2.000 124.455 ;
  RECT 0.000 125.335 2.000 125.395 ;
  RECT 0.000 123.835 2.000 123.955 ;
  RECT 0.000 123.395 2.000 123.455 ;
  RECT 0.000 124.335 2.000 124.395 ;
  RECT 0.000 122.835 2.000 122.955 ;
  RECT 0.000 122.395 2.000 122.455 ;
  RECT 0.000 123.335 2.000 123.395 ;
  RECT 0.000 121.835 2.000 121.955 ;
  RECT 0.000 121.395 2.000 121.455 ;
  RECT 0.000 122.335 2.000 122.395 ;
  RECT 0.000 120.835 2.000 120.955 ;
  RECT 0.000 120.395 2.000 120.455 ;
  RECT 0.000 121.335 2.000 121.395 ;
  RECT 0.000 119.835 2.000 119.955 ;
  RECT 0.000 119.395 2.000 119.455 ;
  RECT 0.000 120.335 2.000 120.395 ;
  RECT 0.000 118.835 2.000 118.955 ;
  RECT 0.000 118.395 2.000 118.455 ;
  RECT 0.000 119.335 2.000 119.395 ;
  RECT 0.000 117.835 2.000 117.955 ;
  RECT 0.000 117.395 2.000 117.455 ;
  RECT 0.000 118.335 2.000 118.395 ;
  RECT 0.000 116.835 2.000 116.955 ;
  RECT 0.000 116.395 2.000 116.455 ;
  RECT 0.000 117.335 2.000 117.395 ;
  RECT 0.000 115.835 2.000 115.955 ;
  RECT 0.000 115.395 2.000 115.455 ;
  RECT 0.000 116.335 2.000 116.395 ;
  RECT 0.000 114.835 2.000 114.955 ;
  RECT 0.000 114.395 2.000 114.455 ;
  RECT 0.000 115.335 2.000 115.395 ;
  RECT 0.000 113.835 2.000 113.955 ;
  RECT 0.000 113.395 2.000 113.455 ;
  RECT 0.000 114.335 2.000 114.395 ;
  RECT 0.000 112.835 2.000 112.955 ;
  RECT 0.000 112.395 2.000 112.455 ;
  RECT 0.000 113.335 2.000 113.395 ;
  RECT 0.000 111.835 2.000 111.955 ;
  RECT 0.000 111.395 2.000 111.455 ;
  RECT 0.000 112.335 2.000 112.395 ;
  RECT 0.000 110.835 2.000 110.955 ;
  RECT 0.000 110.395 2.000 110.455 ;
  RECT 0.000 111.335 2.000 111.395 ;
  RECT 0.000 109.835 2.000 109.955 ;
  RECT 0.000 109.395 2.000 109.455 ;
  RECT 0.000 110.335 2.000 110.395 ;
  RECT 0.000 108.835 2.000 108.955 ;
  RECT 0.000 108.395 2.000 108.455 ;
  RECT 0.000 109.335 2.000 109.395 ;
  RECT 0.000 107.835 2.000 107.955 ;
  RECT 0.000 107.395 2.000 107.455 ;
  RECT 0.000 108.335 2.000 108.395 ;
  RECT 0.000 106.835 2.000 106.955 ;
  RECT 0.000 106.395 2.000 106.455 ;
  RECT 0.000 107.335 2.000 107.395 ;
  RECT 0.000 105.835 2.000 105.955 ;
  RECT 0.000 105.395 2.000 105.455 ;
  RECT 0.000 106.335 2.000 106.395 ;
  RECT 0.000 104.835 2.000 104.955 ;
  RECT 0.000 104.395 2.000 104.455 ;
  RECT 0.000 105.335 2.000 105.395 ;
  RECT 0.000 103.835 2.000 103.955 ;
  RECT 0.000 103.395 2.000 103.455 ;
  RECT 0.000 104.335 2.000 104.395 ;
  RECT 0.000 102.835 2.000 102.955 ;
  RECT 0.000 102.395 2.000 102.455 ;
  RECT 0.000 103.335 2.000 103.395 ;
  RECT 0.000 101.835 2.000 101.955 ;
  RECT 0.000 101.395 2.000 101.455 ;
  RECT 0.000 102.335 2.000 102.395 ;
  RECT 0.000 100.835 2.000 100.955 ;
  RECT 0.000 100.395 2.000 100.455 ;
  RECT 0.000 101.335 2.000 101.395 ;
  RECT 0.000 99.835 2.000 99.955 ;
  RECT 0.000 99.395 2.000 99.455 ;
  RECT 0.000 100.335 2.000 100.395 ;
  RECT 0.000 98.835 2.000 98.955 ;
  RECT 0.000 98.395 2.000 98.455 ;
  RECT 0.000 99.335 2.000 99.395 ;
  RECT 0.000 97.835 2.000 97.955 ;
  RECT 0.000 97.395 2.000 97.455 ;
  RECT 0.000 98.335 2.000 98.395 ;
  RECT 0.000 96.835 2.000 96.955 ;
  RECT 0.000 96.395 2.000 96.455 ;
  RECT 0.000 97.335 2.000 97.395 ;
  RECT 0.000 95.835 2.000 95.955 ;
  RECT 0.000 95.395 2.000 95.455 ;
  RECT 0.000 96.335 2.000 96.395 ;
  RECT 0.000 94.835 2.000 94.955 ;
  RECT 0.000 94.395 2.000 94.455 ;
  RECT 0.000 95.335 2.000 95.395 ;
  RECT 0.000 94.325 2.000 94.395 ;
  RECT 0.000 93.595 2.000 93.665 ;
  RECT 0.000 93.795 2.000 93.935 ;
  RECT 0.000 93.035 2.000 93.155 ;
  RECT 0.000 92.595 2.000 92.655 ;
  RECT 0.000 93.535 2.000 93.595 ;
  RECT 0.000 92.035 2.000 92.155 ;
  RECT 0.000 91.595 2.000 91.655 ;
  RECT 0.000 92.535 2.000 92.595 ;
  RECT 0.000 91.035 2.000 91.155 ;
  RECT 0.000 90.595 2.000 90.655 ;
  RECT 0.000 91.535 2.000 91.595 ;
  RECT 0.000 90.035 2.000 90.155 ;
  RECT 0.000 89.595 2.000 89.655 ;
  RECT 0.000 90.535 2.000 90.595 ;
  RECT 0.000 89.035 2.000 89.155 ;
  RECT 0.000 88.595 2.000 88.655 ;
  RECT 0.000 89.535 2.000 89.595 ;
  RECT 0.000 88.035 2.000 88.155 ;
  RECT 0.000 87.595 2.000 87.655 ;
  RECT 0.000 88.535 2.000 88.595 ;
  RECT 0.000 87.035 2.000 87.155 ;
  RECT 0.000 86.595 2.000 86.655 ;
  RECT 0.000 87.535 2.000 87.595 ;
  RECT 0.000 86.035 2.000 86.155 ;
  RECT 0.000 85.595 2.000 85.655 ;
  RECT 0.000 86.535 2.000 86.595 ;
  RECT 0.000 85.035 2.000 85.155 ;
  RECT 0.000 84.595 2.000 84.655 ;
  RECT 0.000 85.535 2.000 85.595 ;
  RECT 0.000 84.035 2.000 84.155 ;
  RECT 0.000 83.595 2.000 83.655 ;
  RECT 0.000 84.535 2.000 84.595 ;
  RECT 0.000 83.035 2.000 83.155 ;
  RECT 0.000 82.595 2.000 82.655 ;
  RECT 0.000 83.535 2.000 83.595 ;
  RECT 0.000 82.035 2.000 82.155 ;
  RECT 0.000 81.595 2.000 81.655 ;
  RECT 0.000 82.535 2.000 82.595 ;
  RECT 0.000 81.035 2.000 81.155 ;
  RECT 0.000 80.595 2.000 80.655 ;
  RECT 0.000 81.535 2.000 81.595 ;
  RECT 0.000 80.035 2.000 80.155 ;
  RECT 0.000 79.595 2.000 79.655 ;
  RECT 0.000 80.535 2.000 80.595 ;
  RECT 0.000 79.035 2.000 79.155 ;
  RECT 0.000 78.595 2.000 78.655 ;
  RECT 0.000 79.535 2.000 79.595 ;
  RECT 0.000 78.035 2.000 78.155 ;
  RECT 0.000 77.595 2.000 77.655 ;
  RECT 0.000 78.535 2.000 78.595 ;
  RECT 0.000 77.035 2.000 77.155 ;
  RECT 0.000 76.595 2.000 76.655 ;
  RECT 0.000 77.535 2.000 77.595 ;
  RECT 0.000 76.035 2.000 76.155 ;
  RECT 0.000 75.595 2.000 75.655 ;
  RECT 0.000 76.535 2.000 76.595 ;
  RECT 0.000 75.035 2.000 75.155 ;
  RECT 0.000 74.595 2.000 74.655 ;
  RECT 0.000 75.535 2.000 75.595 ;
  RECT 0.000 74.035 2.000 74.155 ;
  RECT 0.000 73.595 2.000 73.655 ;
  RECT 0.000 74.535 2.000 74.595 ;
  RECT 0.000 73.035 2.000 73.155 ;
  RECT 0.000 72.595 2.000 72.655 ;
  RECT 0.000 73.535 2.000 73.595 ;
  RECT 0.000 72.035 2.000 72.155 ;
  RECT 0.000 71.595 2.000 71.655 ;
  RECT 0.000 72.535 2.000 72.595 ;
  RECT 0.000 71.035 2.000 71.155 ;
  RECT 0.000 70.595 2.000 70.655 ;
  RECT 0.000 71.535 2.000 71.595 ;
  RECT 0.000 70.035 2.000 70.155 ;
  RECT 0.000 69.595 2.000 69.655 ;
  RECT 0.000 70.535 2.000 70.595 ;
  RECT 0.000 69.035 2.000 69.155 ;
  RECT 0.000 68.595 2.000 68.655 ;
  RECT 0.000 69.535 2.000 69.595 ;
  RECT 0.000 68.035 2.000 68.155 ;
  RECT 0.000 67.595 2.000 67.655 ;
  RECT 0.000 68.535 2.000 68.595 ;
  RECT 0.000 67.035 2.000 67.155 ;
  RECT 0.000 66.595 2.000 66.655 ;
  RECT 0.000 67.535 2.000 67.595 ;
  RECT 0.000 66.035 2.000 66.155 ;
  RECT 0.000 65.595 2.000 65.655 ;
  RECT 0.000 66.535 2.000 66.595 ;
  RECT 0.000 65.035 2.000 65.155 ;
  RECT 0.000 64.595 2.000 64.655 ;
  RECT 0.000 65.535 2.000 65.595 ;
  RECT 0.000 64.035 2.000 64.155 ;
  RECT 0.000 63.595 2.000 63.655 ;
  RECT 0.000 64.535 2.000 64.595 ;
  RECT 0.000 63.035 2.000 63.155 ;
  RECT 0.000 62.595 2.000 62.655 ;
  RECT 0.000 63.535 2.000 63.595 ;
  RECT 0.000 62.035 2.000 62.155 ;
  RECT 0.000 61.595 2.000 61.655 ;
  RECT 0.000 62.535 2.000 62.595 ;
  RECT 0.000 61.525 2.000 61.595 ;
  RECT 0.000 60.795 2.000 60.865 ;
  RECT 0.000 60.995 2.000 61.135 ;
  RECT 0.000 60.235 2.000 60.355 ;
  RECT 0.000 59.795 2.000 59.855 ;
  RECT 0.000 60.735 2.000 60.795 ;
  RECT 0.000 59.235 2.000 59.355 ;
  RECT 0.000 58.795 2.000 58.855 ;
  RECT 0.000 59.735 2.000 59.795 ;
  RECT 0.000 58.235 2.000 58.355 ;
  RECT 0.000 57.795 2.000 57.855 ;
  RECT 0.000 58.735 2.000 58.795 ;
  RECT 0.000 57.235 2.000 57.355 ;
  RECT 0.000 56.795 2.000 56.855 ;
  RECT 0.000 57.735 2.000 57.795 ;
  RECT 0.000 56.235 2.000 56.355 ;
  RECT 0.000 55.795 2.000 55.855 ;
  RECT 0.000 56.735 2.000 56.795 ;
  RECT 0.000 55.235 2.000 55.355 ;
  RECT 0.000 54.795 2.000 54.855 ;
  RECT 0.000 55.735 2.000 55.795 ;
  RECT 0.000 54.235 2.000 54.355 ;
  RECT 0.000 53.795 2.000 53.855 ;
  RECT 0.000 54.735 2.000 54.795 ;
  RECT 0.000 53.235 2.000 53.355 ;
  RECT 0.000 52.795 2.000 52.855 ;
  RECT 0.000 53.735 2.000 53.795 ;
  RECT 0.000 52.235 2.000 52.355 ;
  RECT 0.000 51.795 2.000 51.855 ;
  RECT 0.000 52.735 2.000 52.795 ;
  RECT 0.000 51.235 2.000 51.355 ;
  RECT 0.000 50.795 2.000 50.855 ;
  RECT 0.000 51.735 2.000 51.795 ;
  RECT 0.000 50.235 2.000 50.355 ;
  RECT 0.000 49.795 2.000 49.855 ;
  RECT 0.000 50.735 2.000 50.795 ;
  RECT 0.000 49.235 2.000 49.355 ;
  RECT 0.000 48.795 2.000 48.855 ;
  RECT 0.000 49.735 2.000 49.795 ;
  RECT 0.000 48.235 2.000 48.355 ;
  RECT 0.000 47.795 2.000 47.855 ;
  RECT 0.000 48.735 2.000 48.795 ;
  RECT 0.000 47.235 2.000 47.355 ;
  RECT 0.000 46.795 2.000 46.855 ;
  RECT 0.000 47.735 2.000 47.795 ;
  RECT 0.000 46.235 2.000 46.355 ;
  RECT 0.000 45.795 2.000 45.855 ;
  RECT 0.000 46.735 2.000 46.795 ;
  RECT 0.000 45.235 2.000 45.355 ;
  RECT 0.000 44.795 2.000 44.855 ;
  RECT 0.000 45.735 2.000 45.795 ;
  RECT 0.000 44.235 2.000 44.355 ;
  RECT 0.000 43.795 2.000 43.855 ;
  RECT 0.000 44.735 2.000 44.795 ;
  RECT 0.000 43.235 2.000 43.355 ;
  RECT 0.000 42.795 2.000 42.855 ;
  RECT 0.000 43.735 2.000 43.795 ;
  RECT 0.000 42.235 2.000 42.355 ;
  RECT 0.000 41.795 2.000 41.855 ;
  RECT 0.000 42.735 2.000 42.795 ;
  RECT 0.000 41.235 2.000 41.355 ;
  RECT 0.000 40.795 2.000 40.855 ;
  RECT 0.000 41.735 2.000 41.795 ;
  RECT 0.000 40.235 2.000 40.355 ;
  RECT 0.000 39.795 2.000 39.855 ;
  RECT 0.000 40.735 2.000 40.795 ;
  RECT 0.000 39.235 2.000 39.355 ;
  RECT 0.000 38.795 2.000 38.855 ;
  RECT 0.000 39.735 2.000 39.795 ;
  RECT 0.000 38.235 2.000 38.355 ;
  RECT 0.000 37.795 2.000 37.855 ;
  RECT 0.000 38.735 2.000 38.795 ;
  RECT 0.000 37.235 2.000 37.355 ;
  RECT 0.000 36.795 2.000 36.855 ;
  RECT 0.000 37.735 2.000 37.795 ;
  RECT 0.000 36.235 2.000 36.355 ;
  RECT 0.000 35.795 2.000 35.855 ;
  RECT 0.000 36.735 2.000 36.795 ;
  RECT 0.000 35.235 2.000 35.355 ;
  RECT 0.000 34.795 2.000 34.855 ;
  RECT 0.000 35.735 2.000 35.795 ;
  RECT 0.000 34.235 2.000 34.355 ;
  RECT 0.000 33.795 2.000 33.855 ;
  RECT 0.000 34.735 2.000 34.795 ;
  RECT 0.000 33.235 2.000 33.355 ;
  RECT 0.000 32.795 2.000 32.855 ;
  RECT 0.000 33.735 2.000 33.795 ;
  RECT 0.000 32.235 2.000 32.355 ;
  RECT 0.000 31.795 2.000 31.855 ;
  RECT 0.000 32.735 2.000 32.795 ;
  RECT 0.000 31.235 2.000 31.355 ;
  RECT 0.000 30.795 2.000 30.855 ;
  RECT 0.000 31.735 2.000 31.795 ;
  RECT 0.000 30.235 2.000 30.355 ;
  RECT 0.000 29.795 2.000 29.855 ;
  RECT 0.000 30.735 2.000 30.795 ;
  RECT 0.000 29.235 2.000 29.355 ;
  RECT 0.000 28.795 2.000 28.855 ;
  RECT 0.000 29.735 2.000 29.795 ;
  RECT 0.000 28.715 2.000 28.795 ;
  RECT 0.000 28.195 2.000 28.335 ;
END
END SYLA55_512X32X4CM2
END LIBRARY






