//======================================================
// Copyright (C) 2020 By 
// All Rights Reserved
//======================================================
// Module : 
// Author : 
// Contact : 
// Date : 
//=======================================================
// Description :
//========================================================
`ifndef DEFINE
  `define DEFINE
  
// `define DATA_WIDTH 8
// `define ADDR_WIDTH 8
// `define FLAG_WIDTH 32
// `define PORT_WIDTH 128
`define TOT_DATA   40959
`define TOT_FLAG   10239

`endif
